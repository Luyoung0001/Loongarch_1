module WallaceTree32x32 (
    input clk,
    input reset,
    input mult,
    input  [31:0] pp0,  pp1,  pp2,  pp3,  pp4,  pp5,  pp6,  pp7,
                   pp8,  pp9,  pp10, pp11, pp12, pp13, pp14, pp15,
                   pp16, pp17, pp18, pp19, pp20, pp21, pp22, pp23,
                   pp24, pp25, pp26, pp27, pp28, pp29, pp30, pp31,
    output reg [63:0] opa,
    output reg [63:0] opb,
    output reg done
);
 wire	[31: 0]	Fir1_S, Fir1_C;
 wire	[31: 0]	Fir2_S, Fir2_C;
 wire	[31: 0]	Fir3_S, Fir3_C;
 wire	[31: 0]	Fir4_S, Fir4_C;
 wire	[31: 0]	Fir5_S, Fir5_C;
 wire	[31: 0]	Fir6_S, Fir6_C;
 wire	[31: 0]	Fir7_S, Fir7_C;
 wire	[31: 0]	Fir8_S, Fir8_C;
 wire	[31: 0]	Fir9_S, Fir9_C;
 wire	[31: 0]	Fir10_S, Fir10_C;
 wire	[30: 0]	Fir11_S, Fir11_C;

  HalfAdder fir1ha0 ( pp0[1], pp1[0], Fir1_S[0], Fir1_C[0] );
  FullAdder  fir1fa1 ( pp0[2],   pp1[1],    pp2[0],
                       Fir1_S[1],   Fir1_C[1] );
  FullAdder fir1fa2  ( pp0[3],    pp1[2],    pp2[1],
                      Fir1_S[2],   Fir1_C[2] );
  FullAdder fir1fa3  ( pp0[4],    pp1[3],    pp2[2],
                      Fir1_S[3],   Fir1_C[3] );
  FullAdder fir1fa4  ( pp0[5],    pp1[4],    pp2[3],
                      Fir1_S[4],   Fir1_C[4] );
  FullAdder fir1fa5  ( pp0[6],    pp1[5],    pp2[4],
                      Fir1_S[5],   Fir1_C[5] );
  FullAdder fir1fa6  ( pp0[7],    pp1[6],    pp2[5],
                      Fir1_S[6],   Fir1_C[6] );
  FullAdder fir1fa7  ( pp0[8],    pp1[7],    pp2[6],
                      Fir1_S[7],   Fir1_C[7] );
  FullAdder fir1fa8  ( pp0[9],    pp1[8],    pp2[7],
                      Fir1_S[8],   Fir1_C[8] );
  FullAdder fir1fa9  ( pp0[10],    pp1[9],    pp2[8],
                      Fir1_S[9],   Fir1_C[9] );
  FullAdder fir1fa10 ( pp0[11],   pp1[10],    pp2[9],
                      Fir1_S[10],  Fir1_C[10] );
  FullAdder fir1fa11 ( pp0[12],   pp1[11],   pp2[10],
                      Fir1_S[11],  Fir1_C[11] );
  FullAdder fir1fa12 ( pp0[13],   pp1[12],   pp2[11],
                      Fir1_S[12],  Fir1_C[12] );
  FullAdder fir1fa13 ( pp0[14],   pp1[13],   pp2[12],
                      Fir1_S[13],  Fir1_C[13] );
  FullAdder fir1fa14 ( pp0[15],   pp1[14],   pp2[13],
                      Fir1_S[14],  Fir1_C[14] );
  FullAdder fir1fa15 ( pp0[16],   pp1[15],   pp2[14],
                      Fir1_S[15],  Fir1_C[15] );
  FullAdder fir1fa16 ( pp0[17],   pp1[16],   pp2[15],
                      Fir1_S[16],  Fir1_C[16] );
  FullAdder fir1fa17 ( pp0[18],   pp1[17],   pp2[16],
                      Fir1_S[17],  Fir1_C[17] );
  FullAdder fir1fa18 ( pp0[19],   pp1[18],   pp2[17],
                      Fir1_S[18],  Fir1_C[18] );
  FullAdder fir1fa19 ( pp0[20],   pp1[19],   pp2[18],
                      Fir1_S[19],  Fir1_C[19] );
  FullAdder fir1fa20 ( pp0[21],   pp1[20],   pp2[19],
                      Fir1_S[20],  Fir1_C[20] );
  FullAdder fir1fa21 ( pp0[22],   pp1[21],   pp2[20],
                      Fir1_S[21],  Fir1_C[21] );
  FullAdder fir1fa22 ( pp0[23],   pp1[22],   pp2[21],
                      Fir1_S[22],  Fir1_C[22] );
  FullAdder fir1fa23 ( pp0[24],   pp1[23],   pp2[22],
                      Fir1_S[23],  Fir1_C[23] );
  FullAdder fir1fa24 ( pp0[25],   pp1[24],   pp2[23],
                      Fir1_S[24],  Fir1_C[24] );
  FullAdder fir1fa25 ( pp0[26],   pp1[25],   pp2[24],
                      Fir1_S[25],  Fir1_C[25] );
  FullAdder fir1fa26 ( pp0[27],   pp1[26],   pp2[25],
                      Fir1_S[26],  Fir1_C[26] );
  FullAdder fir1fa27 ( pp0[28],   pp1[27],   pp2[26],
                      Fir1_S[27],  Fir1_C[27] );
  FullAdder fir1fa28 ( pp0[29],   pp1[28],   pp2[27],
                      Fir1_S[28],  Fir1_C[28] );
  FullAdder fir1fa29 ( pp0[30],   pp1[29],   pp2[28],
                      Fir1_S[29],  Fir1_C[29] );
  FullAdder fir1fa30 ( pp0[31],   pp1[30],   pp2[29],
                      Fir1_S[30],  Fir1_C[30] );
  HalfAdder fir1ha31 ( pp1[31],   pp2[30],
                      Fir1_S[31],  Fir1_C[31] );

HalfAdder fir2ha0 ( pp3[1], pp4[0], Fir2_S[0], Fir2_C[0] );
  FullAdder  fir2fa1 ( pp3[2],   pp4[1],    pp5[0],
                       Fir2_S[1],   Fir2_C[1] );
  FullAdder fir2fa2  ( pp3[3],    pp4[2],    pp5[1],
                      Fir2_S[2],   Fir2_C[2] );
  FullAdder fir2fa3  ( pp3[4],    pp4[3],    pp5[2],
                      Fir2_S[3],   Fir2_C[3] );
  FullAdder fir2fa4  ( pp3[5],    pp4[4],    pp5[3],
                      Fir2_S[4],   Fir2_C[4] );
  FullAdder fir2fa5  ( pp3[6],    pp4[5],    pp5[4],
                      Fir2_S[5],   Fir2_C[5] );
  FullAdder fir2fa6  ( pp3[7],    pp4[6],    pp5[5],
                      Fir2_S[6],   Fir2_C[6] );
  FullAdder fir2fa7  ( pp3[8],    pp4[7],    pp5[6],
                      Fir2_S[7],   Fir2_C[7] );
  FullAdder fir2fa8  ( pp3[9],    pp4[8],    pp5[7],
                      Fir2_S[8],   Fir2_C[8] );
  FullAdder fir2fa9  ( pp3[10],    pp4[9],    pp5[8],
                      Fir2_S[9],   Fir2_C[9] );
  FullAdder fir2fa10 ( pp3[11],   pp4[10],    pp5[9],
                      Fir2_S[10],  Fir2_C[10] );
  FullAdder fir2fa11 ( pp3[12],   pp4[11],   pp5[10],
                      Fir2_S[11],  Fir2_C[11] );
  FullAdder fir2fa12 ( pp3[13],   pp4[12],   pp5[11],
                      Fir2_S[12],  Fir2_C[12] );
  FullAdder fir2fa13 ( pp3[14],   pp4[13],   pp5[12],
                      Fir2_S[13],  Fir2_C[13] );
  FullAdder fir2fa14 ( pp3[15],   pp4[14],   pp5[13],
                      Fir2_S[14],  Fir2_C[14] );
  FullAdder fir2fa15 ( pp3[16],   pp4[15],   pp5[14],
                      Fir2_S[15],  Fir2_C[15] );
  FullAdder fir2fa16 ( pp3[17],   pp4[16],   pp5[15],
                      Fir2_S[16],  Fir2_C[16] );
  FullAdder fir2fa17 ( pp3[18],   pp4[17],   pp5[16],
                      Fir2_S[17],  Fir2_C[17] );
  FullAdder fir2fa18 ( pp3[19],   pp4[18],   pp5[17],
                      Fir2_S[18],  Fir2_C[18] );
  FullAdder fir2fa19 ( pp3[20],   pp4[19],   pp5[18],
                      Fir2_S[19],  Fir2_C[19] );
  FullAdder fir2fa20 ( pp3[21],   pp4[20],   pp5[19],
                      Fir2_S[20],  Fir2_C[20] );
  FullAdder fir2fa21 ( pp3[22],   pp4[21],   pp5[20],
                      Fir2_S[21],  Fir2_C[21] );
  FullAdder fir2fa22 ( pp3[23],   pp4[22],   pp5[21],
                      Fir2_S[22],  Fir2_C[22] );
  FullAdder fir2fa23 ( pp3[24],   pp4[23],   pp5[22],
                      Fir2_S[23],  Fir2_C[23] );
  FullAdder fir2fa24 ( pp3[25],   pp4[24],   pp5[23],
                      Fir2_S[24],  Fir2_C[24] );
  FullAdder fir2fa25 ( pp3[26],   pp4[25],   pp5[24],
                      Fir2_S[25],  Fir2_C[25] );
  FullAdder fir2fa26 ( pp3[27],   pp4[26],   pp5[25],
                      Fir2_S[26],  Fir2_C[26] );
  FullAdder fir2fa27 ( pp3[28],   pp4[27],   pp5[26],
                      Fir2_S[27],  Fir2_C[27] );
  FullAdder fir2fa28 ( pp3[29],   pp4[28],   pp5[27],
                      Fir2_S[28],  Fir2_C[28] );
  FullAdder fir2fa29 ( pp3[30],   pp4[29],   pp5[28],
                      Fir2_S[29],  Fir2_C[29] );
  FullAdder fir2fa30 ( pp3[31],   pp4[30],   pp5[29],
                      Fir2_S[30],  Fir2_C[30] );
  HalfAdder fir2ha31 ( pp4[31],   pp5[30],
                      Fir2_S[31],  Fir2_C[31] );

HalfAdder fir3ha0 ( pp6[1], pp7[0], Fir3_S[0], Fir3_C[0] );
  FullAdder  fir3fa1 ( pp6[2],   pp7[1],    pp8[0],
                       Fir3_S[1],   Fir3_C[1] );
  FullAdder fir3fa2  ( pp6[3],    pp7[2],    pp8[1],
                      Fir3_S[2],   Fir3_C[2] );
  FullAdder fir3fa3  ( pp6[4],    pp7[3],    pp8[2],
                      Fir3_S[3],   Fir3_C[3] );
  FullAdder fir3fa4  ( pp6[5],    pp7[4],    pp8[3],
                      Fir3_S[4],   Fir3_C[4] );
  FullAdder fir3fa5  ( pp6[6],    pp7[5],    pp8[4],
                      Fir3_S[5],   Fir3_C[5] );
  FullAdder fir3fa6  ( pp6[7],    pp7[6],    pp8[5],
                      Fir3_S[6],   Fir3_C[6] );
  FullAdder fir3fa7  ( pp6[8],    pp7[7],    pp8[6],
                      Fir3_S[7],   Fir3_C[7] );
  FullAdder fir3fa8  ( pp6[9],    pp7[8],    pp8[7],
                      Fir3_S[8],   Fir3_C[8] );
  FullAdder fir3fa9  ( pp6[10],    pp7[9],    pp8[8],
                      Fir3_S[9],   Fir3_C[9] );
  FullAdder fir3fa10 ( pp6[11],   pp7[10],    pp8[9],
                      Fir3_S[10],  Fir3_C[10] );
  FullAdder fir3fa11 ( pp6[12],   pp7[11],   pp8[10],
                      Fir3_S[11],  Fir3_C[11] );
  FullAdder fir3fa12 ( pp6[13],   pp7[12],   pp8[11],
                      Fir3_S[12],  Fir3_C[12] );
  FullAdder fir3fa13 ( pp6[14],   pp7[13],   pp8[12],
                      Fir3_S[13],  Fir3_C[13] );
  FullAdder fir3fa14 ( pp6[15],   pp7[14],   pp8[13],
                      Fir3_S[14],  Fir3_C[14] );
  FullAdder fir3fa15 ( pp6[16],   pp7[15],   pp8[14],
                      Fir3_S[15],  Fir3_C[15] );
  FullAdder fir3fa16 ( pp6[17],   pp7[16],   pp8[15],
                      Fir3_S[16],  Fir3_C[16] );
  FullAdder fir3fa17 ( pp6[18],   pp7[17],   pp8[16],
                      Fir3_S[17],  Fir3_C[17] );
  FullAdder fir3fa18 ( pp6[19],   pp7[18],   pp8[17],
                      Fir3_S[18],  Fir3_C[18] );
  FullAdder fir3fa19 ( pp6[20],   pp7[19],   pp8[18],
                      Fir3_S[19],  Fir3_C[19] );
  FullAdder fir3fa20 ( pp6[21],   pp7[20],   pp8[19],
                      Fir3_S[20],  Fir3_C[20] );
  FullAdder fir3fa21 ( pp6[22],   pp7[21],   pp8[20],
                      Fir3_S[21],  Fir3_C[21] );
  FullAdder fir3fa22 ( pp6[23],   pp7[22],   pp8[21],
                      Fir3_S[22],  Fir3_C[22] );
  FullAdder fir3fa23 ( pp6[24],   pp7[23],   pp8[22],
                      Fir3_S[23],  Fir3_C[23] );
  FullAdder fir3fa24 ( pp6[25],   pp7[24],   pp8[23],
                      Fir3_S[24],  Fir3_C[24] );
  FullAdder fir3fa25 ( pp6[26],   pp7[25],   pp8[24],
                      Fir3_S[25],  Fir3_C[25] );
  FullAdder fir3fa26 ( pp6[27],   pp7[26],   pp8[25],
                      Fir3_S[26],  Fir3_C[26] );
  FullAdder fir3fa27 ( pp6[28],   pp7[27],   pp8[26],
                      Fir3_S[27],  Fir3_C[27] );
  FullAdder fir3fa28 ( pp6[29],   pp7[28],   pp8[27],
                      Fir3_S[28],  Fir3_C[28] );
  FullAdder fir3fa29 ( pp6[30],   pp7[29],   pp8[28],
                      Fir3_S[29],  Fir3_C[29] );
  FullAdder fir3fa30 ( pp6[31],   pp7[30],   pp8[29],
                      Fir3_S[30],  Fir3_C[30] );
  HalfAdder fir3ha31 ( pp7[31],   pp8[30],
                      Fir3_S[31],  Fir3_C[31] );

HalfAdder fir4ha0 ( pp9[1], pp10[0], Fir4_S[0], Fir4_C[0] );
  FullAdder  fir4fa1 ( pp9[2],   pp10[1],    pp11[0],
                       Fir4_S[1],   Fir4_C[1] );
  FullAdder fir4fa2  ( pp9[3],    pp10[2],    pp11[1],
                      Fir4_S[2],   Fir4_C[2] );
  FullAdder fir4fa3  ( pp9[4],    pp10[3],    pp11[2],
                      Fir4_S[3],   Fir4_C[3] );
  FullAdder fir4fa4  ( pp9[5],    pp10[4],    pp11[3],
                      Fir4_S[4],   Fir4_C[4] );
  FullAdder fir4fa5  ( pp9[6],    pp10[5],    pp11[4],
                      Fir4_S[5],   Fir4_C[5] );
  FullAdder fir4fa6  ( pp9[7],    pp10[6],    pp11[5],
                      Fir4_S[6],   Fir4_C[6] );
  FullAdder fir4fa7  ( pp9[8],    pp10[7],    pp11[6],
                      Fir4_S[7],   Fir4_C[7] );
  FullAdder fir4fa8  ( pp9[9],    pp10[8],    pp11[7],
                      Fir4_S[8],   Fir4_C[8] );
  FullAdder fir4fa9  ( pp9[10],    pp10[9],    pp11[8],
                      Fir4_S[9],   Fir4_C[9] );
  FullAdder fir4fa10 ( pp9[11],   pp10[10],    pp11[9],
                      Fir4_S[10],  Fir4_C[10] );
  FullAdder fir4fa11 ( pp9[12],   pp10[11],   pp11[10],
                      Fir4_S[11],  Fir4_C[11] );
  FullAdder fir4fa12 ( pp9[13],   pp10[12],   pp11[11],
                      Fir4_S[12],  Fir4_C[12] );
  FullAdder fir4fa13 ( pp9[14],   pp10[13],   pp11[12],
                      Fir4_S[13],  Fir4_C[13] );
  FullAdder fir4fa14 ( pp9[15],   pp10[14],   pp11[13],
                      Fir4_S[14],  Fir4_C[14] );
  FullAdder fir4fa15 ( pp9[16],   pp10[15],   pp11[14],
                      Fir4_S[15],  Fir4_C[15] );
  FullAdder fir4fa16 ( pp9[17],   pp10[16],   pp11[15],
                      Fir4_S[16],  Fir4_C[16] );
  FullAdder fir4fa17 ( pp9[18],   pp10[17],   pp11[16],
                      Fir4_S[17],  Fir4_C[17] );
  FullAdder fir4fa18 ( pp9[19],   pp10[18],   pp11[17],
                      Fir4_S[18],  Fir4_C[18] );
  FullAdder fir4fa19 ( pp9[20],   pp10[19],   pp11[18],
                      Fir4_S[19],  Fir4_C[19] );
  FullAdder fir4fa20 ( pp9[21],   pp10[20],   pp11[19],
                      Fir4_S[20],  Fir4_C[20] );
  FullAdder fir4fa21 ( pp9[22],   pp10[21],   pp11[20],
                      Fir4_S[21],  Fir4_C[21] );
  FullAdder fir4fa22 ( pp9[23],   pp10[22],   pp11[21],
                      Fir4_S[22],  Fir4_C[22] );
  FullAdder fir4fa23 ( pp9[24],   pp10[23],   pp11[22],
                      Fir4_S[23],  Fir4_C[23] );
  FullAdder fir4fa24 ( pp9[25],   pp10[24],   pp11[23],
                      Fir4_S[24],  Fir4_C[24] );
  FullAdder fir4fa25 ( pp9[26],   pp10[25],   pp11[24],
                      Fir4_S[25],  Fir4_C[25] );
  FullAdder fir4fa26 ( pp9[27],   pp10[26],   pp11[25],
                      Fir4_S[26],  Fir4_C[26] );
  FullAdder fir4fa27 ( pp9[28],   pp10[27],   pp11[26],
                      Fir4_S[27],  Fir4_C[27] );
  FullAdder fir4fa28 ( pp9[29],   pp10[28],   pp11[27],
                      Fir4_S[28],  Fir4_C[28] );
  FullAdder fir4fa29 ( pp9[30],   pp10[29],   pp11[28],
                      Fir4_S[29],  Fir4_C[29] );
  FullAdder fir4fa30 ( pp9[31],   pp10[30],   pp11[29],
                      Fir4_S[30],  Fir4_C[30] );
  HalfAdder fir4ha31 ( pp10[31],   pp11[30],
                      Fir4_S[31],  Fir4_C[31] );

HalfAdder fir5ha0 ( pp12[1], pp13[0], Fir5_S[0], Fir5_C[0] );
  FullAdder  fir5fa1 ( pp12[2],   pp13[1],    pp14[0],
                       Fir5_S[1],   Fir5_C[1] );
  FullAdder fir5fa2  ( pp12[3],    pp13[2],    pp14[1],
                      Fir5_S[2],   Fir5_C[2] );
  FullAdder fir5fa3  ( pp12[4],    pp13[3],    pp14[2],
                      Fir5_S[3],   Fir5_C[3] );
  FullAdder fir5fa4  ( pp12[5],    pp13[4],    pp14[3],
                      Fir5_S[4],   Fir5_C[4] );
  FullAdder fir5fa5  ( pp12[6],    pp13[5],    pp14[4],
                      Fir5_S[5],   Fir5_C[5] );
  FullAdder fir5fa6  ( pp12[7],    pp13[6],    pp14[5],
                      Fir5_S[6],   Fir5_C[6] );
  FullAdder fir5fa7  ( pp12[8],    pp13[7],    pp14[6],
                      Fir5_S[7],   Fir5_C[7] );
  FullAdder fir5fa8  ( pp12[9],    pp13[8],    pp14[7],
                      Fir5_S[8],   Fir5_C[8] );
  FullAdder fir5fa9  ( pp12[10],    pp13[9],    pp14[8],
                      Fir5_S[9],   Fir5_C[9] );
  FullAdder fir5fa10 ( pp12[11],   pp13[10],    pp14[9],
                      Fir5_S[10],  Fir5_C[10] );
  FullAdder fir5fa11 ( pp12[12],   pp13[11],   pp14[10],
                      Fir5_S[11],  Fir5_C[11] );
  FullAdder fir5fa12 ( pp12[13],   pp13[12],   pp14[11],
                      Fir5_S[12],  Fir5_C[12] );
  FullAdder fir5fa13 ( pp12[14],   pp13[13],   pp14[12],
                      Fir5_S[13],  Fir5_C[13] );
  FullAdder fir5fa14 ( pp12[15],   pp13[14],   pp14[13],
                      Fir5_S[14],  Fir5_C[14] );
  FullAdder fir5fa15 ( pp12[16],   pp13[15],   pp14[14],
                      Fir5_S[15],  Fir5_C[15] );
  FullAdder fir5fa16 ( pp12[17],   pp13[16],   pp14[15],
                      Fir5_S[16],  Fir5_C[16] );
  FullAdder fir5fa17 ( pp12[18],   pp13[17],   pp14[16],
                      Fir5_S[17],  Fir5_C[17] );
  FullAdder fir5fa18 ( pp12[19],   pp13[18],   pp14[17],
                      Fir5_S[18],  Fir5_C[18] );
  FullAdder fir5fa19 ( pp12[20],   pp13[19],   pp14[18],
                      Fir5_S[19],  Fir5_C[19] );
  FullAdder fir5fa20 ( pp12[21],   pp13[20],   pp14[19],
                      Fir5_S[20],  Fir5_C[20] );
  FullAdder fir5fa21 ( pp12[22],   pp13[21],   pp14[20],
                      Fir5_S[21],  Fir5_C[21] );
  FullAdder fir5fa22 ( pp12[23],   pp13[22],   pp14[21],
                      Fir5_S[22],  Fir5_C[22] );
  FullAdder fir5fa23 ( pp12[24],   pp13[23],   pp14[22],
                      Fir5_S[23],  Fir5_C[23] );
  FullAdder fir5fa24 ( pp12[25],   pp13[24],   pp14[23],
                      Fir5_S[24],  Fir5_C[24] );
  FullAdder fir5fa25 ( pp12[26],   pp13[25],   pp14[24],
                      Fir5_S[25],  Fir5_C[25] );
  FullAdder fir5fa26 ( pp12[27],   pp13[26],   pp14[25],
                      Fir5_S[26],  Fir5_C[26] );
  FullAdder fir5fa27 ( pp12[28],   pp13[27],   pp14[26],
                      Fir5_S[27],  Fir5_C[27] );
  FullAdder fir5fa28 ( pp12[29],   pp13[28],   pp14[27],
                      Fir5_S[28],  Fir5_C[28] );
  FullAdder fir5fa29 ( pp12[30],   pp13[29],   pp14[28],
                      Fir5_S[29],  Fir5_C[29] );
  FullAdder fir5fa30 ( pp12[31],   pp13[30],   pp14[29],
                      Fir5_S[30],  Fir5_C[30] );
  HalfAdder fir5ha31 ( pp13[31],   pp14[30],
                      Fir5_S[31],  Fir5_C[31] );


  HalfAdder fir6ha0 ( pp15[1], pp16[0], Fir6_S[0], Fir6_C[0] );
  FullAdder  fir6fa1 ( pp15[2],   pp16[1],    pp17[0],
                       Fir6_S[1],   Fir6_C[1] );
  FullAdder fir6fa2  ( pp15[3],    pp16[2],    pp17[1],
                      Fir6_S[2],   Fir6_C[2] );
  FullAdder fir6fa3  ( pp15[4],    pp16[3],    pp17[2],
                      Fir6_S[3],   Fir6_C[3] );
  FullAdder fir6fa4  ( pp15[5],    pp16[4],    pp17[3],
                      Fir6_S[4],   Fir6_C[4] );
  FullAdder fir6fa5  ( pp15[6],    pp16[5],    pp17[4],
                      Fir6_S[5],   Fir6_C[5] );
  FullAdder fir6fa6  ( pp15[7],    pp16[6],    pp17[5],
                      Fir6_S[6],   Fir6_C[6] );
  FullAdder fir6fa7  ( pp15[8],    pp16[7],    pp17[6],
                      Fir6_S[7],   Fir6_C[7] );
  FullAdder fir6fa8  ( pp15[9],    pp16[8],    pp17[7],
                      Fir6_S[8],   Fir6_C[8] );
  FullAdder fir6fa9  ( pp15[10],    pp16[9],    pp17[8],
                      Fir6_S[9],   Fir6_C[9] );
  FullAdder fir6fa10 ( pp15[11],   pp16[10],    pp17[9],
                      Fir6_S[10],  Fir6_C[10] );
  FullAdder fir6fa11 ( pp15[12],   pp16[11],   pp17[10],
                      Fir6_S[11],  Fir6_C[11] );
  FullAdder fir6fa12 ( pp15[13],   pp16[12],   pp17[11],
                      Fir6_S[12],  Fir6_C[12] );
  FullAdder fir6fa13 ( pp15[14],   pp16[13],   pp17[12],
                      Fir6_S[13],  Fir6_C[13] );
  FullAdder fir6fa14 ( pp15[15],   pp16[14],   pp17[13],
                      Fir6_S[14],  Fir6_C[14] );
  FullAdder fir6fa15 ( pp15[16],   pp16[15],   pp17[14],
                      Fir6_S[15],  Fir6_C[15] );
  FullAdder fir6fa16 ( pp15[17],   pp16[16],   pp17[15],
                      Fir6_S[16],  Fir6_C[16] );
  FullAdder fir6fa17 ( pp15[18],   pp16[17],   pp17[16],
                      Fir6_S[17],  Fir6_C[17] );
  FullAdder fir6fa18 ( pp15[19],   pp16[18],   pp17[17],
                      Fir6_S[18],  Fir6_C[18] );
  FullAdder fir6fa19 ( pp15[20],   pp16[19],   pp17[18],
                      Fir6_S[19],  Fir6_C[19] );
  FullAdder fir6fa20 ( pp15[21],   pp16[20],   pp17[19],
                      Fir6_S[20],  Fir6_C[20] );
  FullAdder fir6fa21 ( pp15[22],   pp16[21],   pp17[20],
                      Fir6_S[21],  Fir6_C[21] );
  FullAdder fir6fa22 ( pp15[23],   pp16[22],   pp17[21],
                      Fir6_S[22],  Fir6_C[22] );
  FullAdder fir6fa23 ( pp15[24],   pp16[23],   pp17[22],
                      Fir6_S[23],  Fir6_C[23] );
  FullAdder fir6fa24 ( pp15[25],   pp16[24],   pp17[23],
                      Fir6_S[24],  Fir6_C[24] );
  FullAdder fir6fa25 ( pp15[26],   pp16[25],   pp17[24],
                      Fir6_S[25],  Fir6_C[25] );
  FullAdder fir6fa26 ( pp15[27],   pp16[26],   pp17[25],
                      Fir6_S[26],  Fir6_C[26] );
  FullAdder fir6fa27 ( pp15[28],   pp16[27],   pp17[26],
                      Fir6_S[27],  Fir6_C[27] );
  FullAdder fir6fa28 ( pp15[29],   pp16[28],   pp17[27],
                      Fir6_S[28],  Fir6_C[28] );
  FullAdder fir6fa29 ( pp15[30],   pp16[29],   pp17[28],
                      Fir6_S[29],  Fir6_C[29] );
  FullAdder fir6fa30 ( pp15[31],   pp16[30],   pp17[29],
                      Fir6_S[30],  Fir6_C[30] );
  HalfAdder fir6ha31 ( pp16[31],   pp17[30],
                      Fir6_S[31],  Fir6_C[31] );

  HalfAdder fir7ha0 ( pp18[1], pp19[0], Fir7_S[0], Fir7_C[0] );
  FullAdder  fir7fa1 ( pp18[2],   pp19[1],    pp20[0],
                       Fir7_S[1],   Fir7_C[1] );
  FullAdder fir7fa2  ( pp18[3],    pp19[2],    pp20[1],
                      Fir7_S[2],   Fir7_C[2] );
  FullAdder fir7fa3  ( pp18[4],    pp19[3],    pp20[2],
                      Fir7_S[3],   Fir7_C[3] );
  FullAdder fir7fa4  ( pp18[5],    pp19[4],    pp20[3],
                      Fir7_S[4],   Fir7_C[4] );
  FullAdder fir7fa5  ( pp18[6],    pp19[5],    pp20[4],
                      Fir7_S[5],   Fir7_C[5] );
  FullAdder fir7fa6  ( pp18[7],    pp19[6],    pp20[5],
                      Fir7_S[6],   Fir7_C[6] );
  FullAdder fir7fa7  ( pp18[8],    pp19[7],    pp20[6],
                      Fir7_S[7],   Fir7_C[7] );
  FullAdder fir7fa8  ( pp18[9],    pp19[8],    pp20[7],
                      Fir7_S[8],   Fir7_C[8] );
  FullAdder fir7fa9  ( pp18[10],    pp19[9],    pp20[8],
                      Fir7_S[9],   Fir7_C[9] );
  FullAdder fir7fa10 ( pp18[11],   pp19[10],    pp20[9],
                      Fir7_S[10],  Fir7_C[10] );
  FullAdder fir7fa11 ( pp18[12],   pp19[11],   pp20[10],
                      Fir7_S[11],  Fir7_C[11] );
  FullAdder fir7fa12 ( pp18[13],   pp19[12],   pp20[11],
                      Fir7_S[12],  Fir7_C[12] );
  FullAdder fir7fa13 ( pp18[14],   pp19[13],   pp20[12],
                      Fir7_S[13],  Fir7_C[13] );
  FullAdder fir7fa14 ( pp18[15],   pp19[14],   pp20[13],
                      Fir7_S[14],  Fir7_C[14] );
  FullAdder fir7fa15 ( pp18[16],   pp19[15],   pp20[14],
                      Fir7_S[15],  Fir7_C[15] );
  FullAdder fir7fa16 ( pp18[17],   pp19[16],   pp20[15],
                      Fir7_S[16],  Fir7_C[16] );
  FullAdder fir7fa17 ( pp18[18],   pp19[17],   pp20[16],
                      Fir7_S[17],  Fir7_C[17] );
  FullAdder fir7fa18 ( pp18[19],   pp19[18],   pp20[17],
                      Fir7_S[18],  Fir7_C[18] );
  FullAdder fir7fa19 ( pp18[20],   pp19[19],   pp20[18],
                      Fir7_S[19],  Fir7_C[19] );
  FullAdder fir7fa20 ( pp18[21],   pp19[20],   pp20[19],
                      Fir7_S[20],  Fir7_C[20] );
  FullAdder fir7fa21 ( pp18[22],   pp19[21],   pp20[20],
                      Fir7_S[21],  Fir7_C[21] );
  FullAdder fir7fa22 ( pp18[23],   pp19[22],   pp20[21],
                      Fir7_S[22],  Fir7_C[22] );
  FullAdder fir7fa23 ( pp18[24],   pp19[23],   pp20[22],
                      Fir7_S[23],  Fir7_C[23] );
  FullAdder fir7fa24 ( pp18[25],   pp19[24],   pp20[23],
                      Fir7_S[24],  Fir7_C[24] );
  FullAdder fir7fa25 ( pp18[26],   pp19[25],   pp20[24],
                      Fir7_S[25],  Fir7_C[25] );
  FullAdder fir7fa26 ( pp18[27],   pp19[26],   pp20[25],
                      Fir7_S[26],  Fir7_C[26] );
  FullAdder fir7fa27 ( pp18[28],   pp19[27],   pp20[26],
                      Fir7_S[27],  Fir7_C[27] );
  FullAdder fir7fa28 ( pp18[29],   pp19[28],   pp20[27],
                      Fir7_S[28],  Fir7_C[28] );
  FullAdder fir7fa29 ( pp18[30],   pp19[29],   pp20[28],
                      Fir7_S[29],  Fir7_C[29] );
  FullAdder fir7fa30 ( pp18[31],   pp19[30],   pp20[29],
                      Fir7_S[30],  Fir7_C[30] );
  HalfAdder fir7ha31 ( pp19[31],   pp20[30],
                      Fir7_S[31],  Fir7_C[31] );


HalfAdder fir8ha0 ( pp21[1], pp22[0], Fir8_S[0], Fir8_C[0] );
  FullAdder  fir8fa1 ( pp21[2],   pp22[1],    pp23[0],
                       Fir8_S[1],   Fir8_C[1] );
  FullAdder fir8fa2  ( pp21[3],    pp22[2],    pp23[1],
                      Fir8_S[2],   Fir8_C[2] );
  FullAdder fir8fa3  ( pp21[4],    pp22[3],    pp23[2],
                      Fir8_S[3],   Fir8_C[3] );
  FullAdder fir8fa4  ( pp21[5],    pp22[4],    pp23[3],
                      Fir8_S[4],   Fir8_C[4] );
  FullAdder fir8fa5  ( pp21[6],    pp22[5],    pp23[4],
                      Fir8_S[5],   Fir8_C[5] );
  FullAdder fir8fa6  ( pp21[7],    pp22[6],    pp23[5],
                      Fir8_S[6],   Fir8_C[6] );
  FullAdder fir8fa7  ( pp21[8],    pp22[7],    pp23[6],
                      Fir8_S[7],   Fir8_C[7] );
  FullAdder fir8fa8  ( pp21[9],    pp22[8],    pp23[7],
                      Fir8_S[8],   Fir8_C[8] );
  FullAdder fir8fa9  ( pp21[10],    pp22[9],    pp23[8],
                      Fir8_S[9],   Fir8_C[9] );
  FullAdder fir8fa10 ( pp21[11],   pp22[10],    pp23[9],
                      Fir8_S[10],  Fir8_C[10] );
  FullAdder fir8fa11 ( pp21[12],   pp22[11],   pp23[10],
                      Fir8_S[11],  Fir8_C[11] );
  FullAdder fir8fa12 ( pp21[13],   pp22[12],   pp23[11],
                      Fir8_S[12],  Fir8_C[12] );
  FullAdder fir8fa13 ( pp21[14],   pp22[13],   pp23[12],
                      Fir8_S[13],  Fir8_C[13] );
  FullAdder fir8fa14 ( pp21[15],   pp22[14],   pp23[13],
                      Fir8_S[14],  Fir8_C[14] );
  FullAdder fir8fa15 ( pp21[16],   pp22[15],   pp23[14],
                      Fir8_S[15],  Fir8_C[15] );
  FullAdder fir8fa16 ( pp21[17],   pp22[16],   pp23[15],
                      Fir8_S[16],  Fir8_C[16] );
  FullAdder fir8fa17 ( pp21[18],   pp22[17],   pp23[16],
                      Fir8_S[17],  Fir8_C[17] );
  FullAdder fir8fa18 ( pp21[19],   pp22[18],   pp23[17],
                      Fir8_S[18],  Fir8_C[18] );
  FullAdder fir8fa19 ( pp21[20],   pp22[19],   pp23[18],
                      Fir8_S[19],  Fir8_C[19] );
  FullAdder fir8fa20 ( pp21[21],   pp22[20],   pp23[19],
                      Fir8_S[20],  Fir8_C[20] );
  FullAdder fir8fa21 ( pp21[22],   pp22[21],   pp23[20],
                      Fir8_S[21],  Fir8_C[21] );
  FullAdder fir8fa22 ( pp21[23],   pp22[22],   pp23[21],
                      Fir8_S[22],  Fir8_C[22] );
  FullAdder fir8fa23 ( pp21[24],   pp22[23],   pp23[22],
                      Fir8_S[23],  Fir8_C[23] );
  FullAdder fir8fa24 ( pp21[25],   pp22[24],   pp23[23],
                      Fir8_S[24],  Fir8_C[24] );
  FullAdder fir8fa25 ( pp21[26],   pp22[25],   pp23[24],
                      Fir8_S[25],  Fir8_C[25] );
  FullAdder fir8fa26 ( pp21[27],   pp22[26],   pp23[25],
                      Fir8_S[26],  Fir8_C[26] );
  FullAdder fir8fa27 ( pp21[28],   pp22[27],   pp23[26],
                      Fir8_S[27],  Fir8_C[27] );
  FullAdder fir8fa28 ( pp21[29],   pp22[28],   pp23[27],
                      Fir8_S[28],  Fir8_C[28] );
  FullAdder fir8fa29 ( pp21[30],   pp22[29],   pp23[28],
                      Fir8_S[29],  Fir8_C[29] );
  FullAdder fir8fa30 ( pp21[31],   pp22[30],   pp23[29],
                      Fir8_S[30],  Fir8_C[30] );
  HalfAdder fir8ha31 ( pp22[31],   pp23[30],
                      Fir8_S[31],  Fir8_C[31] );


HalfAdder fir9ha0 ( pp24[1], pp25[0], Fir9_S[0], Fir9_C[0] );
  FullAdder  fir9fa1 ( pp24[2],   pp25[1],    pp26[0],
                       Fir9_S[1],   Fir9_C[1] );
  FullAdder fir9fa2  ( pp24[3],    pp25[2],    pp26[1],
                      Fir9_S[2],   Fir9_C[2] );
  FullAdder fir9fa3  ( pp24[4],    pp25[3],    pp26[2],
                      Fir9_S[3],   Fir9_C[3] );
  FullAdder fir9fa4  ( pp24[5],    pp25[4],    pp26[3],
                      Fir9_S[4],   Fir9_C[4] );
  FullAdder fir9fa5  ( pp24[6],    pp25[5],    pp26[4],
                      Fir9_S[5],   Fir9_C[5] );
  FullAdder fir9fa6  ( pp24[7],    pp25[6],    pp26[5],
                      Fir9_S[6],   Fir9_C[6] );
  FullAdder fir9fa7  ( pp24[8],    pp25[7],    pp26[6],
                      Fir9_S[7],   Fir9_C[7] );
  FullAdder fir9fa8  ( pp24[9],    pp25[8],    pp26[7],
                      Fir9_S[8],   Fir9_C[8] );
  FullAdder fir9fa9  ( pp24[10],    pp25[9],    pp26[8],
                      Fir9_S[9],   Fir9_C[9] );
  FullAdder fir9fa10 ( pp24[11],   pp25[10],    pp26[9],
                      Fir9_S[10],  Fir9_C[10] );
  FullAdder fir9fa11 ( pp24[12],   pp25[11],   pp26[10],
                      Fir9_S[11],  Fir9_C[11] );
  FullAdder fir9fa12 ( pp24[13],   pp25[12],   pp26[11],
                      Fir9_S[12],  Fir9_C[12] );
  FullAdder fir9fa13 ( pp24[14],   pp25[13],   pp26[12],
                      Fir9_S[13],  Fir9_C[13] );
  FullAdder fir9fa14 ( pp24[15],   pp25[14],   pp26[13],
                      Fir9_S[14],  Fir9_C[14] );
  FullAdder fir9fa15 ( pp24[16],   pp25[15],   pp26[14],
                      Fir9_S[15],  Fir9_C[15] );
  FullAdder fir9fa16 ( pp24[17],   pp25[16],   pp26[15],
                      Fir9_S[16],  Fir9_C[16] );
  FullAdder fir9fa17 ( pp24[18],   pp25[17],   pp26[16],
                      Fir9_S[17],  Fir9_C[17] );
  FullAdder fir9fa18 ( pp24[19],   pp25[18],   pp26[17],
                      Fir9_S[18],  Fir9_C[18] );
  FullAdder fir9fa19 ( pp24[20],   pp25[19],   pp26[18],
                      Fir9_S[19],  Fir9_C[19] );
  FullAdder fir9fa20 ( pp24[21],   pp25[20],   pp26[19],
                      Fir9_S[20],  Fir9_C[20] );
  FullAdder fir9fa21 ( pp24[22],   pp25[21],   pp26[20],
                      Fir9_S[21],  Fir9_C[21] );
  FullAdder fir9fa22 ( pp24[23],   pp25[22],   pp26[21],
                      Fir9_S[22],  Fir9_C[22] );
  FullAdder fir9fa23 ( pp24[24],   pp25[23],   pp26[22],
                      Fir9_S[23],  Fir9_C[23] );
  FullAdder fir9fa24 ( pp24[25],   pp25[24],   pp26[23],
                      Fir9_S[24],  Fir9_C[24] );
  FullAdder fir9fa25 ( pp24[26],   pp25[25],   pp26[24],
                      Fir9_S[25],  Fir9_C[25] );
  FullAdder fir9fa26 ( pp24[27],   pp25[26],   pp26[25],
                      Fir9_S[26],  Fir9_C[26] );
  FullAdder fir9fa27 ( pp24[28],   pp25[27],   pp26[26],
                      Fir9_S[27],  Fir9_C[27] );
  FullAdder fir9fa28 ( pp24[29],   pp25[28],   pp26[27],
                      Fir9_S[28],  Fir9_C[28] );
  FullAdder fir9fa29 ( pp24[30],   pp25[29],   pp26[28],
                      Fir9_S[29],  Fir9_C[29] );
  FullAdder fir9fa30 ( pp24[31],   pp25[30],   pp26[29],
                      Fir9_S[30],  Fir9_C[30] );
  HalfAdder fir9ha31 ( pp25[31],   pp26[30],
                      Fir9_S[31],  Fir9_C[31] );


HalfAdder fir10ha0 ( pp27[1], pp28[0], Fir10_S[0], Fir10_C[0] );
  FullAdder  fir10fa1 ( pp27[2],   pp28[1],    pp29[0],
                       Fir10_S[1],   Fir10_C[1] );
  FullAdder fir10fa2  ( pp27[3],    pp28[2],    pp29[1],
                      Fir10_S[2],   Fir10_C[2] );
  FullAdder fir10fa3  ( pp27[4],    pp28[3],    pp29[2],
                      Fir10_S[3],   Fir10_C[3] );
  FullAdder fir10fa4  ( pp27[5],    pp28[4],    pp29[3],
                      Fir10_S[4],   Fir10_C[4] );
  FullAdder fir10fa5  ( pp27[6],    pp28[5],    pp29[4],
                      Fir10_S[5],   Fir10_C[5] );
  FullAdder fir10fa6  ( pp27[7],    pp28[6],    pp29[5],
                      Fir10_S[6],   Fir10_C[6] );
  FullAdder fir10fa7  ( pp27[8],    pp28[7],    pp29[6],
                      Fir10_S[7],   Fir10_C[7] );
  FullAdder fir10fa8  ( pp27[9],    pp28[8],    pp29[7],
                      Fir10_S[8],   Fir10_C[8] );
  FullAdder fir10fa9  ( pp27[10],    pp28[9],    pp29[8],
                      Fir10_S[9],   Fir10_C[9] );
  FullAdder fir10fa10 ( pp27[11],   pp28[10],    pp29[9],
                      Fir10_S[10],  Fir10_C[10] );
  FullAdder fir10fa11 ( pp27[12],   pp28[11],   pp29[10],
                      Fir10_S[11],  Fir10_C[11] );
  FullAdder fir10fa12 ( pp27[13],   pp28[12],   pp29[11],
                      Fir10_S[12],  Fir10_C[12] );
  FullAdder fir10fa13 ( pp27[14],   pp28[13],   pp29[12],
                      Fir10_S[13],  Fir10_C[13] );
  FullAdder fir10fa14 ( pp27[15],   pp28[14],   pp29[13],
                      Fir10_S[14],  Fir10_C[14] );
  FullAdder fir10fa15 ( pp27[16],   pp28[15],   pp29[14],
                      Fir10_S[15],  Fir10_C[15] );
  FullAdder fir10fa16 ( pp27[17],   pp28[16],   pp29[15],
                      Fir10_S[16],  Fir10_C[16] );
  FullAdder fir10fa17 ( pp27[18],   pp28[17],   pp29[16],
                      Fir10_S[17],  Fir10_C[17] );
  FullAdder fir10fa18 ( pp27[19],   pp28[18],   pp29[17],
                      Fir10_S[18],  Fir10_C[18] );
  FullAdder fir10fa19 ( pp27[20],   pp28[19],   pp29[18],
                      Fir10_S[19],  Fir10_C[19] );
  FullAdder fir10fa20 ( pp27[21],   pp28[20],   pp29[19],
                      Fir10_S[20],  Fir10_C[20] );
  FullAdder fir10fa21 ( pp27[22],   pp28[21],   pp29[20],
                      Fir10_S[21],  Fir10_C[21] );
  FullAdder fir10fa22 ( pp27[23],   pp28[22],   pp29[21],
                      Fir10_S[22],  Fir10_C[22] );
  FullAdder fir10fa23 ( pp27[24],   pp28[23],   pp29[22],
                      Fir10_S[23],  Fir10_C[23] );
  FullAdder fir10fa24 ( pp27[25],   pp28[24],   pp29[23],
                      Fir10_S[24],  Fir10_C[24] );
  FullAdder fir10fa25 ( pp27[26],   pp28[25],   pp29[24],
                      Fir10_S[25],  Fir10_C[25] );
  FullAdder fir10fa26 ( pp27[27],   pp28[26],   pp29[25],
                      Fir10_S[26],  Fir10_C[26] );
  FullAdder fir10fa27 ( pp27[28],   pp28[27],   pp29[26],
                      Fir10_S[27],  Fir10_C[27] );
  FullAdder fir10fa28 ( pp27[29],   pp28[28],   pp29[27],
                      Fir10_S[28],  Fir10_C[28] );
  FullAdder fir10fa29 ( pp27[30],   pp28[29],   pp29[28],
                      Fir10_S[29],  Fir10_C[29] );
  FullAdder fir10fa30 ( pp27[31],   pp28[30],   pp29[29],
                      Fir10_S[30],  Fir10_C[30] );
  HalfAdder fir10ha31 ( pp28[31],   pp29[30],
                      Fir10_S[31],  Fir10_C[31] );

HalfAdder fir11ha0 ( pp30[1], pp31[0], Fir11_S[0], Fir11_C[0] );
HalfAdder fir11ha1 ( pp30[2], pp31[1], Fir11_S[1], Fir11_C[1] );
HalfAdder fir11ha2 ( pp30[3], pp31[2], Fir11_S[2], Fir11_C[2] );
HalfAdder fir11ha3 ( pp30[4], pp31[3], Fir11_S[3], Fir11_C[3] );
HalfAdder fir11ha4 ( pp30[5], pp31[4], Fir11_S[4], Fir11_C[4] );
HalfAdder fir11ha5 ( pp30[6], pp31[5], Fir11_S[5], Fir11_C[5] );
HalfAdder fir11ha6 ( pp30[7], pp31[6], Fir11_S[6], Fir11_C[6] );
HalfAdder fir11ha7 ( pp30[8], pp31[7], Fir11_S[7], Fir11_C[7] );
HalfAdder fir11ha8 ( pp30[9], pp31[8], Fir11_S[8], Fir11_C[8] );
HalfAdder fir11ha9 ( pp30[10], pp31[9], Fir11_S[9], Fir11_C[9] );
HalfAdder fir11ha10 ( pp30[11], pp31[10], Fir11_S[10], Fir11_C[10] );
HalfAdder fir11ha11 ( pp30[12], pp31[11], Fir11_S[11], Fir11_C[11] );
HalfAdder fir11ha12 ( pp30[13], pp31[12], Fir11_S[12], Fir11_C[12] );
HalfAdder fir11ha13 ( pp30[14], pp31[13], Fir11_S[13], Fir11_C[13] );
HalfAdder fir11ha14 ( pp30[15], pp31[14], Fir11_S[14], Fir11_C[14] );
HalfAdder fir11ha15 ( pp30[16], pp31[15], Fir11_S[15], Fir11_C[15] );
HalfAdder fir11ha16 ( pp30[17], pp31[16], Fir11_S[16], Fir11_C[16] );
HalfAdder fir11ha17 ( pp30[18], pp31[17], Fir11_S[17], Fir11_C[17] );
HalfAdder fir11ha18 ( pp30[19], pp31[18], Fir11_S[18], Fir11_C[18] );
HalfAdder fir11ha19 ( pp30[20], pp31[19], Fir11_S[19], Fir11_C[19] );
HalfAdder fir11ha20 ( pp30[21], pp31[20], Fir11_S[20], Fir11_C[20] );
HalfAdder fir11ha21 ( pp30[22], pp31[21], Fir11_S[21], Fir11_C[21] );
HalfAdder fir11ha22 ( pp30[23], pp31[22], Fir11_S[22], Fir11_C[22] );
HalfAdder fir11ha23 ( pp30[24], pp31[23], Fir11_S[23], Fir11_C[23] );
HalfAdder fir11ha24 ( pp30[25], pp31[24], Fir11_S[24], Fir11_C[24] );
HalfAdder fir11ha25 ( pp30[26], pp31[25], Fir11_S[25], Fir11_C[25] );
HalfAdder fir11ha26 ( pp30[27], pp31[26], Fir11_S[26], Fir11_C[26] );
HalfAdder fir11ha27 ( pp30[28], pp31[27], Fir11_S[27], Fir11_C[27] );
HalfAdder fir11ha28 ( pp30[29], pp31[28], Fir11_S[28], Fir11_C[28] );
HalfAdder fir11ha29 ( pp30[30], pp31[29], Fir11_S[29], Fir11_C[29] );
HalfAdder fir11ha30 ( pp30[31], pp31[30], Fir11_S[30], Fir11_C[30] );



 reg	[31: 0]	Fir1_S_, Fir1_C_;
 reg	[31: 0]	Fir2_S_, Fir2_C_;
 reg	[31: 0]	Fir3_S_, Fir3_C_;
 reg	[31: 0]	Fir4_S_, Fir4_C_;
 reg	[31: 0]	Fir5_S_, Fir5_C_;
 reg	[31: 0]	Fir6_S_, Fir6_C_;
 reg	[31: 0]	Fir7_S_, Fir7_C_;
 reg	[31: 0]	Fir8_S_, Fir8_C_;
 reg	[31: 0]	Fir9_S_, Fir9_C_;
 reg	[31: 0]	Fir10_S_, Fir10_C_;
 reg	[30: 0]	Fir11_S_, Fir11_C_;
reg done0;
reg state_done0;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Fir1_S_  <= 32'b0; Fir1_C_  <= 32'b0;
        Fir2_S_  <= 32'b0; Fir2_C_  <= 32'b0;
        Fir3_S_  <= 32'b0; Fir3_C_  <= 32'b0;
        Fir4_S_  <= 32'b0; Fir4_C_  <= 32'b0;
        Fir5_S_  <= 32'b0; Fir5_C_  <= 32'b0;
        Fir6_S_  <= 32'b0; Fir6_C_  <= 32'b0;
        Fir7_S_  <= 32'b0; Fir7_C_  <= 32'b0;
        Fir8_S_  <= 32'b0; Fir8_C_  <= 32'b0;
        Fir9_S_  <= 32'b0; Fir9_C_  <= 32'b0;
        Fir10_S_ <= 32'b0; Fir10_C_ <= 32'b0;
        Fir11_S_ <= 31'b0; Fir11_C_ <= 31'b0;
        done0    <= 1'b0;
        state_done0 <= 1'b0;
    end else begin
        case (state_done0)
            1'b0: begin
                if (mult) begin
                    Fir1_S_  <= Fir1_S;   Fir1_C_  <= Fir1_C;
                    Fir2_S_  <= Fir2_S;   Fir2_C_  <= Fir2_C;
                    Fir3_S_  <= Fir3_S;   Fir3_C_  <= Fir3_C;
                    Fir4_S_  <= Fir4_S;   Fir4_C_  <= Fir4_C;
                    Fir5_S_  <= Fir5_S;   Fir5_C_  <= Fir5_C;
                    Fir6_S_  <= Fir6_S;   Fir6_C_  <= Fir6_C;
                    Fir7_S_  <= Fir7_S;   Fir7_C_  <= Fir7_C;
                    Fir8_S_  <= Fir8_S;   Fir8_C_  <= Fir8_C;
                    Fir9_S_  <= Fir9_S;   Fir9_C_  <= Fir9_C;
                    Fir10_S_ <= Fir10_S;  Fir10_C_ <= Fir10_C;
                    Fir11_S_ <= Fir11_S;  Fir11_C_ <= Fir11_C;
                    done0 <= 1'b1;
                    state_done0 <= 1'b1;
                end else begin
                    done0 <= 1'b0;
                end
            end
            1'b1: begin
                done0 <= 1'b0; 
                if (!mult) begin
                    state_done0 <= 1'b0;
                end
            end
        endcase
    end
end


  //===================Second stage===============================

wire	[31: 0]	Sec1_S_, Sec1_C_;
wire	[31: 0]	Sec2_S_, Sec2_C_;
wire	[31: 0]	Sec3_S_, Sec3_C_;
wire	[31: 0]	Sec4_S_, Sec4_C_;
wire	[31: 0]	Sec5_S_, Sec5_C_;
wire	[31: 0]	Sec6_S_, Sec6_C_;
wire	[31: 0]	Sec7_S_, Sec7_C_;
wire	[31: 0]	Sec8_S_, Sec8_C_;
wire	[31: 0]	Sec9_S_, Sec9_C_;
wire	[31: 0]	Sec10_S_, Sec10_C_;
wire	[30: 0]	Sec11_S_, Sec11_C_;


HalfAdder sec1ha0( Fir1_S_[1], Fir1_C_[0], Sec1_S_[0], Sec1_C_[0] );
HalfAdder sec1ha1( Fir1_S_[2], Fir1_C_[1], Sec1_S_[1], Sec1_C_[1] );
HalfAdder sec1ha2( Fir1_S_[3], Fir1_C_[2], Sec1_S_[2], Sec1_C_[2] );
HalfAdder sec1ha3( Fir1_S_[4], Fir1_C_[3], Sec1_S_[3], Sec1_C_[3] );
HalfAdder sec1ha4( Fir1_S_[5], Fir1_C_[4], Sec1_S_[4], Sec1_C_[4] );
HalfAdder sec1ha5( Fir1_S_[6], Fir1_C_[5], Sec1_S_[5], Sec1_C_[5] );
HalfAdder sec1ha6( Fir1_S_[7], Fir1_C_[6], Sec1_S_[6], Sec1_C_[6] );
HalfAdder sec1ha7( Fir1_S_[8], Fir1_C_[7], Sec1_S_[7], Sec1_C_[7] );
HalfAdder sec1ha8( Fir1_S_[9], Fir1_C_[8], Sec1_S_[8], Sec1_C_[8] );
HalfAdder sec1ha9( Fir1_S_[10], Fir1_C_[9], Sec1_S_[9], Sec1_C_[9] );
HalfAdder sec1ha10( Fir1_S_[11], Fir1_C_[10], Sec1_S_[10], Sec1_C_[10] );
HalfAdder sec1ha11( Fir1_S_[12], Fir1_C_[11], Sec1_S_[11], Sec1_C_[11] );
HalfAdder sec1ha12( Fir1_S_[13], Fir1_C_[12], Sec1_S_[12], Sec1_C_[12] );
HalfAdder sec1ha13( Fir1_S_[14], Fir1_C_[13], Sec1_S_[13], Sec1_C_[13] );
HalfAdder sec1ha14( Fir1_S_[15], Fir1_C_[14], Sec1_S_[14], Sec1_C_[14] );
HalfAdder sec1ha15( Fir1_S_[16], Fir1_C_[15], Sec1_S_[15], Sec1_C_[15] );
HalfAdder sec1ha16( Fir1_S_[17], Fir1_C_[16], Sec1_S_[16], Sec1_C_[16] );
HalfAdder sec1ha17( Fir1_S_[18], Fir1_C_[17], Sec1_S_[17], Sec1_C_[17] );
HalfAdder sec1ha18( Fir1_S_[19], Fir1_C_[18], Sec1_S_[18], Sec1_C_[18] );
HalfAdder sec1ha19( Fir1_S_[20], Fir1_C_[19], Sec1_S_[19], Sec1_C_[19] );
HalfAdder sec1ha20( Fir1_S_[21], Fir1_C_[20], Sec1_S_[20], Sec1_C_[20] );
HalfAdder sec1ha21( Fir1_S_[22], Fir1_C_[21], Sec1_S_[21], Sec1_C_[21] );
HalfAdder sec1ha22( Fir1_S_[23], Fir1_C_[22], Sec1_S_[22], Sec1_C_[22] );
HalfAdder sec1ha23( Fir1_S_[24], Fir1_C_[23], Sec1_S_[23], Sec1_C_[23] );
HalfAdder sec1ha24( Fir1_S_[25], Fir1_C_[24], Sec1_S_[24], Sec1_C_[24] );
HalfAdder sec1ha25( Fir1_S_[26], Fir1_C_[25], Sec1_S_[25], Sec1_C_[25] );
HalfAdder sec1ha26( Fir1_S_[27], Fir1_C_[26], Sec1_S_[26], Sec1_C_[26] );
HalfAdder sec1ha27( Fir1_S_[28], Fir1_C_[27], Sec1_S_[27], Sec1_C_[27] );
HalfAdder sec1ha28( Fir1_S_[29], Fir1_C_[28], Sec1_S_[28], Sec1_C_[28] );
HalfAdder sec1ha29( Fir1_S_[30], Fir1_C_[29], Sec1_S_[29], Sec1_C_[29] );
HalfAdder sec1ha30( Fir1_S_[31], Fir1_C_[30], Sec1_S_[30], Sec1_C_[30] );
HalfAdder sec1ha31( pp2[31], Fir1_C_[31], Sec1_S_[31], Sec1_C_[31] );

HalfAdder sec2ha0( Fir2_S_[1], Fir2_C_[0], Sec2_S_[0], Sec2_C_[0] );
HalfAdder sec2ha1( Fir2_S_[2], Fir2_C_[1], Sec2_S_[1], Sec2_C_[1] );
HalfAdder sec2ha2( Fir2_S_[3], Fir2_C_[2], Sec2_S_[2], Sec2_C_[2] );
HalfAdder sec2ha3( Fir2_S_[4], Fir2_C_[3], Sec2_S_[3], Sec2_C_[3] );
HalfAdder sec2ha4( Fir2_S_[5], Fir2_C_[4], Sec2_S_[4], Sec2_C_[4] );
HalfAdder sec2ha5( Fir2_S_[6], Fir2_C_[5], Sec2_S_[5], Sec2_C_[5] );
HalfAdder sec2ha6( Fir2_S_[7], Fir2_C_[6], Sec2_S_[6], Sec2_C_[6] );
HalfAdder sec2ha7( Fir2_S_[8], Fir2_C_[7], Sec2_S_[7], Sec2_C_[7] );
HalfAdder sec2ha8( Fir2_S_[9], Fir2_C_[8], Sec2_S_[8], Sec2_C_[8] );
HalfAdder sec2ha9( Fir2_S_[10], Fir2_C_[9], Sec2_S_[9], Sec2_C_[9] );
HalfAdder sec2ha10( Fir2_S_[11], Fir2_C_[10], Sec2_S_[10], Sec2_C_[10] );
HalfAdder sec2ha11( Fir2_S_[12], Fir2_C_[11], Sec2_S_[11], Sec2_C_[11] );
HalfAdder sec2ha12( Fir2_S_[13], Fir2_C_[12], Sec2_S_[12], Sec2_C_[12] );
HalfAdder sec2ha13( Fir2_S_[14], Fir2_C_[13], Sec2_S_[13], Sec2_C_[13] );
HalfAdder sec2ha14( Fir2_S_[15], Fir2_C_[14], Sec2_S_[14], Sec2_C_[14] );
HalfAdder sec2ha15( Fir2_S_[16], Fir2_C_[15], Sec2_S_[15], Sec2_C_[15] );
HalfAdder sec2ha16( Fir2_S_[17], Fir2_C_[16], Sec2_S_[16], Sec2_C_[16] );
HalfAdder sec2ha17( Fir2_S_[18], Fir2_C_[17], Sec2_S_[17], Sec2_C_[17] );
HalfAdder sec2ha18( Fir2_S_[19], Fir2_C_[18], Sec2_S_[18], Sec2_C_[18] );
HalfAdder sec2ha19( Fir2_S_[20], Fir2_C_[19], Sec2_S_[19], Sec2_C_[19] );
HalfAdder sec2ha20( Fir2_S_[21], Fir2_C_[20], Sec2_S_[20], Sec2_C_[20] );
HalfAdder sec2ha21( Fir2_S_[22], Fir2_C_[21], Sec2_S_[21], Sec2_C_[21] );
HalfAdder sec2ha22( Fir2_S_[23], Fir2_C_[22], Sec2_S_[22], Sec2_C_[22] );
HalfAdder sec2ha23( Fir2_S_[24], Fir2_C_[23], Sec2_S_[23], Sec2_C_[23] );
HalfAdder sec2ha24( Fir2_S_[25], Fir2_C_[24], Sec2_S_[24], Sec2_C_[24] );
HalfAdder sec2ha25( Fir2_S_[26], Fir2_C_[25], Sec2_S_[25], Sec2_C_[25] );
HalfAdder sec2ha26( Fir2_S_[27], Fir2_C_[26], Sec2_S_[26], Sec2_C_[26] );
HalfAdder sec2ha27( Fir2_S_[28], Fir2_C_[27], Sec2_S_[27], Sec2_C_[27] );
HalfAdder sec2ha28( Fir2_S_[29], Fir2_C_[28], Sec2_S_[28], Sec2_C_[28] );
HalfAdder sec2ha29( Fir2_S_[30], Fir2_C_[29], Sec2_S_[29], Sec2_C_[29] );
HalfAdder sec2ha30( Fir2_S_[31], Fir2_C_[30], Sec2_S_[30], Sec2_C_[30] );
HalfAdder sec2ha31( pp5[31], Fir2_C_[31], Sec2_S_[31], Sec2_C_[31] );


HalfAdder sec3ha0( Fir3_S_[1], Fir3_C_[0], Sec3_S_[0], Sec3_C_[0] );
HalfAdder sec3ha1( Fir3_S_[2], Fir3_C_[1], Sec3_S_[1], Sec3_C_[1] );
HalfAdder sec3ha2( Fir3_S_[3], Fir3_C_[2], Sec3_S_[2], Sec3_C_[2] );
HalfAdder sec3ha3( Fir3_S_[4], Fir3_C_[3], Sec3_S_[3], Sec3_C_[3] );
HalfAdder sec3ha4( Fir3_S_[5], Fir3_C_[4], Sec3_S_[4], Sec3_C_[4] );
HalfAdder sec3ha5( Fir3_S_[6], Fir3_C_[5], Sec3_S_[5], Sec3_C_[5] );
HalfAdder sec3ha6( Fir3_S_[7], Fir3_C_[6], Sec3_S_[6], Sec3_C_[6] );
HalfAdder sec3ha7( Fir3_S_[8], Fir3_C_[7], Sec3_S_[7], Sec3_C_[7] );
HalfAdder sec3ha8( Fir3_S_[9], Fir3_C_[8], Sec3_S_[8], Sec3_C_[8] );
HalfAdder sec3ha9( Fir3_S_[10], Fir3_C_[9], Sec3_S_[9], Sec3_C_[9] );
HalfAdder sec3ha10( Fir3_S_[11], Fir3_C_[10], Sec3_S_[10], Sec3_C_[10] );
HalfAdder sec3ha11( Fir3_S_[12], Fir3_C_[11], Sec3_S_[11], Sec3_C_[11] );
HalfAdder sec3ha12( Fir3_S_[13], Fir3_C_[12], Sec3_S_[12], Sec3_C_[12] );
HalfAdder sec3ha13( Fir3_S_[14], Fir3_C_[13], Sec3_S_[13], Sec3_C_[13] );
HalfAdder sec3ha14( Fir3_S_[15], Fir3_C_[14], Sec3_S_[14], Sec3_C_[14] );
HalfAdder sec3ha15( Fir3_S_[16], Fir3_C_[15], Sec3_S_[15], Sec3_C_[15] );
HalfAdder sec3ha16( Fir3_S_[17], Fir3_C_[16], Sec3_S_[16], Sec3_C_[16] );
HalfAdder sec3ha17( Fir3_S_[18], Fir3_C_[17], Sec3_S_[17], Sec3_C_[17] );
HalfAdder sec3ha18( Fir3_S_[19], Fir3_C_[18], Sec3_S_[18], Sec3_C_[18] );
HalfAdder sec3ha19( Fir3_S_[20], Fir3_C_[19], Sec3_S_[19], Sec3_C_[19] );
HalfAdder sec3ha20( Fir3_S_[21], Fir3_C_[20], Sec3_S_[20], Sec3_C_[20] );
HalfAdder sec3ha21( Fir3_S_[22], Fir3_C_[21], Sec3_S_[21], Sec3_C_[21] );
HalfAdder sec3ha22( Fir3_S_[23], Fir3_C_[22], Sec3_S_[22], Sec3_C_[22] );
HalfAdder sec3ha23( Fir3_S_[24], Fir3_C_[23], Sec3_S_[23], Sec3_C_[23] );
HalfAdder sec3ha24( Fir3_S_[25], Fir3_C_[24], Sec3_S_[24], Sec3_C_[24] );
HalfAdder sec3ha25( Fir3_S_[26], Fir3_C_[25], Sec3_S_[25], Sec3_C_[25] );
HalfAdder sec3ha26( Fir3_S_[27], Fir3_C_[26], Sec3_S_[26], Sec3_C_[26] );
HalfAdder sec3ha27( Fir3_S_[28], Fir3_C_[27], Sec3_S_[27], Sec3_C_[27] );
HalfAdder sec3ha28( Fir3_S_[29], Fir3_C_[28], Sec3_S_[28], Sec3_C_[28] );
HalfAdder sec3ha29( Fir3_S_[30], Fir3_C_[29], Sec3_S_[29], Sec3_C_[29] );
HalfAdder sec3ha30( Fir3_S_[31], Fir3_C_[30], Sec3_S_[30], Sec3_C_[30] );
HalfAdder sec3ha31( pp8[31], Fir3_C_[31], Sec3_S_[31], Sec3_C_[31] );

HalfAdder sec4ha0( Fir4_S_[1], Fir4_C_[0], Sec4_S_[0], Sec4_C_[0] );
HalfAdder sec4ha1( Fir4_S_[2], Fir4_C_[1], Sec4_S_[1], Sec4_C_[1] );
HalfAdder sec4ha2( Fir4_S_[3], Fir4_C_[2], Sec4_S_[2], Sec4_C_[2] );
HalfAdder sec4ha3( Fir4_S_[4], Fir4_C_[3], Sec4_S_[3], Sec4_C_[3] );
HalfAdder sec4ha4( Fir4_S_[5], Fir4_C_[4], Sec4_S_[4], Sec4_C_[4] );
HalfAdder sec4ha5( Fir4_S_[6], Fir4_C_[5], Sec4_S_[5], Sec4_C_[5] );
HalfAdder sec4ha6( Fir4_S_[7], Fir4_C_[6], Sec4_S_[6], Sec4_C_[6] );
HalfAdder sec4ha7( Fir4_S_[8], Fir4_C_[7], Sec4_S_[7], Sec4_C_[7] );
HalfAdder sec4ha8( Fir4_S_[9], Fir4_C_[8], Sec4_S_[8], Sec4_C_[8] );
HalfAdder sec4ha9( Fir4_S_[10], Fir4_C_[9], Sec4_S_[9], Sec4_C_[9] );
HalfAdder sec4ha10( Fir4_S_[11], Fir4_C_[10], Sec4_S_[10], Sec4_C_[10] );
HalfAdder sec4ha11( Fir4_S_[12], Fir4_C_[11], Sec4_S_[11], Sec4_C_[11] );
HalfAdder sec4ha12( Fir4_S_[13], Fir4_C_[12], Sec4_S_[12], Sec4_C_[12] );
HalfAdder sec4ha13( Fir4_S_[14], Fir4_C_[13], Sec4_S_[13], Sec4_C_[13] );
HalfAdder sec4ha14( Fir4_S_[15], Fir4_C_[14], Sec4_S_[14], Sec4_C_[14] );
HalfAdder sec4ha15( Fir4_S_[16], Fir4_C_[15], Sec4_S_[15], Sec4_C_[15] );
HalfAdder sec4ha16( Fir4_S_[17], Fir4_C_[16], Sec4_S_[16], Sec4_C_[16] );
HalfAdder sec4ha17( Fir4_S_[18], Fir4_C_[17], Sec4_S_[17], Sec4_C_[17] );
HalfAdder sec4ha18( Fir4_S_[19], Fir4_C_[18], Sec4_S_[18], Sec4_C_[18] );
HalfAdder sec4ha19( Fir4_S_[20], Fir4_C_[19], Sec4_S_[19], Sec4_C_[19] );
HalfAdder sec4ha20( Fir4_S_[21], Fir4_C_[20], Sec4_S_[20], Sec4_C_[20] );
HalfAdder sec4ha21( Fir4_S_[22], Fir4_C_[21], Sec4_S_[21], Sec4_C_[21] );
HalfAdder sec4ha22( Fir4_S_[23], Fir4_C_[22], Sec4_S_[22], Sec4_C_[22] );
HalfAdder sec4ha23( Fir4_S_[24], Fir4_C_[23], Sec4_S_[23], Sec4_C_[23] );
HalfAdder sec4ha24( Fir4_S_[25], Fir4_C_[24], Sec4_S_[24], Sec4_C_[24] );
HalfAdder sec4ha25( Fir4_S_[26], Fir4_C_[25], Sec4_S_[25], Sec4_C_[25] );
HalfAdder sec4ha26( Fir4_S_[27], Fir4_C_[26], Sec4_S_[26], Sec4_C_[26] );
HalfAdder sec4ha27( Fir4_S_[28], Fir4_C_[27], Sec4_S_[27], Sec4_C_[27] );
HalfAdder sec4ha28( Fir4_S_[29], Fir4_C_[28], Sec4_S_[28], Sec4_C_[28] );
HalfAdder sec4ha29( Fir4_S_[30], Fir4_C_[29], Sec4_S_[29], Sec4_C_[29] );
HalfAdder sec4ha30( Fir4_S_[31], Fir4_C_[30], Sec4_S_[30], Sec4_C_[30] );
HalfAdder sec4ha31( pp11[31], Fir4_C_[31], Sec4_S_[31], Sec4_C_[31] );


HalfAdder sec5ha0( Fir5_S_[1], Fir5_C_[0], Sec5_S_[0], Sec5_C_[0] );
HalfAdder sec5ha1( Fir5_S_[2], Fir5_C_[1], Sec5_S_[1], Sec5_C_[1] );
HalfAdder sec5ha2( Fir5_S_[3], Fir5_C_[2], Sec5_S_[2], Sec5_C_[2] );
HalfAdder sec5ha3( Fir5_S_[4], Fir5_C_[3], Sec5_S_[3], Sec5_C_[3] );
HalfAdder sec5ha4( Fir5_S_[5], Fir5_C_[4], Sec5_S_[4], Sec5_C_[4] );
HalfAdder sec5ha5( Fir5_S_[6], Fir5_C_[5], Sec5_S_[5], Sec5_C_[5] );
HalfAdder sec5ha6( Fir5_S_[7], Fir5_C_[6], Sec5_S_[6], Sec5_C_[6] );
HalfAdder sec5ha7( Fir5_S_[8], Fir5_C_[7], Sec5_S_[7], Sec5_C_[7] );
HalfAdder sec5ha8( Fir5_S_[9], Fir5_C_[8], Sec5_S_[8], Sec5_C_[8] );
HalfAdder sec5ha9( Fir5_S_[10], Fir5_C_[9], Sec5_S_[9], Sec5_C_[9] );
HalfAdder sec5ha10( Fir5_S_[11], Fir5_C_[10], Sec5_S_[10], Sec5_C_[10] );
HalfAdder sec5ha11( Fir5_S_[12], Fir5_C_[11], Sec5_S_[11], Sec5_C_[11] );
HalfAdder sec5ha12( Fir5_S_[13], Fir5_C_[12], Sec5_S_[12], Sec5_C_[12] );
HalfAdder sec5ha13( Fir5_S_[14], Fir5_C_[13], Sec5_S_[13], Sec5_C_[13] );
HalfAdder sec5ha14( Fir5_S_[15], Fir5_C_[14], Sec5_S_[14], Sec5_C_[14] );
HalfAdder sec5ha15( Fir5_S_[16], Fir5_C_[15], Sec5_S_[15], Sec5_C_[15] );
HalfAdder sec5ha16( Fir5_S_[17], Fir5_C_[16], Sec5_S_[16], Sec5_C_[16] );
HalfAdder sec5ha17( Fir5_S_[18], Fir5_C_[17], Sec5_S_[17], Sec5_C_[17] );
HalfAdder sec5ha18( Fir5_S_[19], Fir5_C_[18], Sec5_S_[18], Sec5_C_[18] );
HalfAdder sec5ha19( Fir5_S_[20], Fir5_C_[19], Sec5_S_[19], Sec5_C_[19] );
HalfAdder sec5ha20( Fir5_S_[21], Fir5_C_[20], Sec5_S_[20], Sec5_C_[20] );
HalfAdder sec5ha21( Fir5_S_[22], Fir5_C_[21], Sec5_S_[21], Sec5_C_[21] );
HalfAdder sec5ha22( Fir5_S_[23], Fir5_C_[22], Sec5_S_[22], Sec5_C_[22] );
HalfAdder sec5ha23( Fir5_S_[24], Fir5_C_[23], Sec5_S_[23], Sec5_C_[23] );
HalfAdder sec5ha24( Fir5_S_[25], Fir5_C_[24], Sec5_S_[24], Sec5_C_[24] );
HalfAdder sec5ha25( Fir5_S_[26], Fir5_C_[25], Sec5_S_[25], Sec5_C_[25] );
HalfAdder sec5ha26( Fir5_S_[27], Fir5_C_[26], Sec5_S_[26], Sec5_C_[26] );
HalfAdder sec5ha27( Fir5_S_[28], Fir5_C_[27], Sec5_S_[27], Sec5_C_[27] );
HalfAdder sec5ha28( Fir5_S_[29], Fir5_C_[28], Sec5_S_[28], Sec5_C_[28] );
HalfAdder sec5ha29( Fir5_S_[30], Fir5_C_[29], Sec5_S_[29], Sec5_C_[29] );
HalfAdder sec5ha30( Fir5_S_[31], Fir5_C_[30], Sec5_S_[30], Sec5_C_[30] );
HalfAdder sec5ha31( pp14[31], Fir5_C_[31], Sec5_S_[31], Sec5_C_[31] );

HalfAdder sec6ha0( Fir6_S_[1], Fir6_C_[0], Sec6_S_[0], Sec6_C_[0] );
HalfAdder sec6ha1( Fir6_S_[2], Fir6_C_[1], Sec6_S_[1], Sec6_C_[1] );
HalfAdder sec6ha2( Fir6_S_[3], Fir6_C_[2], Sec6_S_[2], Sec6_C_[2] );
HalfAdder sec6ha3( Fir6_S_[4], Fir6_C_[3], Sec6_S_[3], Sec6_C_[3] );
HalfAdder sec6ha4( Fir6_S_[5], Fir6_C_[4], Sec6_S_[4], Sec6_C_[4] );
HalfAdder sec6ha5( Fir6_S_[6], Fir6_C_[5], Sec6_S_[5], Sec6_C_[5] );
HalfAdder sec6ha6( Fir6_S_[7], Fir6_C_[6], Sec6_S_[6], Sec6_C_[6] );
HalfAdder sec6ha7( Fir6_S_[8], Fir6_C_[7], Sec6_S_[7], Sec6_C_[7] );
HalfAdder sec6ha8( Fir6_S_[9], Fir6_C_[8], Sec6_S_[8], Sec6_C_[8] );
HalfAdder sec6ha9( Fir6_S_[10], Fir6_C_[9], Sec6_S_[9], Sec6_C_[9] );
HalfAdder sec6ha10( Fir6_S_[11], Fir6_C_[10], Sec6_S_[10], Sec6_C_[10] );
HalfAdder sec6ha11( Fir6_S_[12], Fir6_C_[11], Sec6_S_[11], Sec6_C_[11] );
HalfAdder sec6ha12( Fir6_S_[13], Fir6_C_[12], Sec6_S_[12], Sec6_C_[12] );
HalfAdder sec6ha13( Fir6_S_[14], Fir6_C_[13], Sec6_S_[13], Sec6_C_[13] );
HalfAdder sec6ha14( Fir6_S_[15], Fir6_C_[14], Sec6_S_[14], Sec6_C_[14] );
HalfAdder sec6ha15( Fir6_S_[16], Fir6_C_[15], Sec6_S_[15], Sec6_C_[15] );
HalfAdder sec6ha16( Fir6_S_[17], Fir6_C_[16], Sec6_S_[16], Sec6_C_[16] );
HalfAdder sec6ha17( Fir6_S_[18], Fir6_C_[17], Sec6_S_[17], Sec6_C_[17] );
HalfAdder sec6ha18( Fir6_S_[19], Fir6_C_[18], Sec6_S_[18], Sec6_C_[18] );
HalfAdder sec6ha19( Fir6_S_[20], Fir6_C_[19], Sec6_S_[19], Sec6_C_[19] );
HalfAdder sec6ha20( Fir6_S_[21], Fir6_C_[20], Sec6_S_[20], Sec6_C_[20] );
HalfAdder sec6ha21( Fir6_S_[22], Fir6_C_[21], Sec6_S_[21], Sec6_C_[21] );
HalfAdder sec6ha22( Fir6_S_[23], Fir6_C_[22], Sec6_S_[22], Sec6_C_[22] );
HalfAdder sec6ha23( Fir6_S_[24], Fir6_C_[23], Sec6_S_[23], Sec6_C_[23] );
HalfAdder sec6ha24( Fir6_S_[25], Fir6_C_[24], Sec6_S_[24], Sec6_C_[24] );
HalfAdder sec6ha25( Fir6_S_[26], Fir6_C_[25], Sec6_S_[25], Sec6_C_[25] );
HalfAdder sec6ha26( Fir6_S_[27], Fir6_C_[26], Sec6_S_[26], Sec6_C_[26] );
HalfAdder sec6ha27( Fir6_S_[28], Fir6_C_[27], Sec6_S_[27], Sec6_C_[27] );
HalfAdder sec6ha28( Fir6_S_[29], Fir6_C_[28], Sec6_S_[28], Sec6_C_[28] );
HalfAdder sec6ha29( Fir6_S_[30], Fir6_C_[29], Sec6_S_[29], Sec6_C_[29] );
HalfAdder sec6ha30( Fir6_S_[31], Fir6_C_[30], Sec6_S_[30], Sec6_C_[30] );
HalfAdder sec6ha31( pp17[31], Fir6_C_[31], Sec6_S_[31], Sec6_C_[31] );

HalfAdder sec7ha0( Fir7_S_[1], Fir7_C_[0], Sec7_S_[0], Sec7_C_[0] );
HalfAdder sec7ha1( Fir7_S_[2], Fir7_C_[1], Sec7_S_[1], Sec7_C_[1] );
HalfAdder sec7ha2( Fir7_S_[3], Fir7_C_[2], Sec7_S_[2], Sec7_C_[2] );
HalfAdder sec7ha3( Fir7_S_[4], Fir7_C_[3], Sec7_S_[3], Sec7_C_[3] );
HalfAdder sec7ha4( Fir7_S_[5], Fir7_C_[4], Sec7_S_[4], Sec7_C_[4] );
HalfAdder sec7ha5( Fir7_S_[6], Fir7_C_[5], Sec7_S_[5], Sec7_C_[5] );
HalfAdder sec7ha6( Fir7_S_[7], Fir7_C_[6], Sec7_S_[6], Sec7_C_[6] );
HalfAdder sec7ha7( Fir7_S_[8], Fir7_C_[7], Sec7_S_[7], Sec7_C_[7] );
HalfAdder sec7ha8( Fir7_S_[9], Fir7_C_[8], Sec7_S_[8], Sec7_C_[8] );
HalfAdder sec7ha9( Fir7_S_[10], Fir7_C_[9], Sec7_S_[9], Sec7_C_[9] );
HalfAdder sec7ha10( Fir7_S_[11], Fir7_C_[10], Sec7_S_[10], Sec7_C_[10] );
HalfAdder sec7ha11( Fir7_S_[12], Fir7_C_[11], Sec7_S_[11], Sec7_C_[11] );
HalfAdder sec7ha12( Fir7_S_[13], Fir7_C_[12], Sec7_S_[12], Sec7_C_[12] );
HalfAdder sec7ha13( Fir7_S_[14], Fir7_C_[13], Sec7_S_[13], Sec7_C_[13] );
HalfAdder sec7ha14( Fir7_S_[15], Fir7_C_[14], Sec7_S_[14], Sec7_C_[14] );
HalfAdder sec7ha15( Fir7_S_[16], Fir7_C_[15], Sec7_S_[15], Sec7_C_[15] );
HalfAdder sec7ha16( Fir7_S_[17], Fir7_C_[16], Sec7_S_[16], Sec7_C_[16] );
HalfAdder sec7ha17( Fir7_S_[18], Fir7_C_[17], Sec7_S_[17], Sec7_C_[17] );
HalfAdder sec7ha18( Fir7_S_[19], Fir7_C_[18], Sec7_S_[18], Sec7_C_[18] );
HalfAdder sec7ha19( Fir7_S_[20], Fir7_C_[19], Sec7_S_[19], Sec7_C_[19] );
HalfAdder sec7ha20( Fir7_S_[21], Fir7_C_[20], Sec7_S_[20], Sec7_C_[20] );
HalfAdder sec7ha21( Fir7_S_[22], Fir7_C_[21], Sec7_S_[21], Sec7_C_[21] );
HalfAdder sec7ha22( Fir7_S_[23], Fir7_C_[22], Sec7_S_[22], Sec7_C_[22] );
HalfAdder sec7ha23( Fir7_S_[24], Fir7_C_[23], Sec7_S_[23], Sec7_C_[23] );
HalfAdder sec7ha24( Fir7_S_[25], Fir7_C_[24], Sec7_S_[24], Sec7_C_[24] );
HalfAdder sec7ha25( Fir7_S_[26], Fir7_C_[25], Sec7_S_[25], Sec7_C_[25] );
HalfAdder sec7ha26( Fir7_S_[27], Fir7_C_[26], Sec7_S_[26], Sec7_C_[26] );
HalfAdder sec7ha27( Fir7_S_[28], Fir7_C_[27], Sec7_S_[27], Sec7_C_[27] );
HalfAdder sec7ha28( Fir7_S_[29], Fir7_C_[28], Sec7_S_[28], Sec7_C_[28] );
HalfAdder sec7ha29( Fir7_S_[30], Fir7_C_[29], Sec7_S_[29], Sec7_C_[29] );
HalfAdder sec7ha30( Fir7_S_[31], Fir7_C_[30], Sec7_S_[30], Sec7_C_[30] );
HalfAdder sec7ha31( pp20[31], Fir7_C_[31], Sec7_S_[31], Sec7_C_[31] );


HalfAdder sec8ha0( Fir8_S_[1], Fir8_C_[0], Sec8_S_[0], Sec8_C_[0] );
HalfAdder sec8ha1( Fir8_S_[2], Fir8_C_[1], Sec8_S_[1], Sec8_C_[1] );
HalfAdder sec8ha2( Fir8_S_[3], Fir8_C_[2], Sec8_S_[2], Sec8_C_[2] );
HalfAdder sec8ha3( Fir8_S_[4], Fir8_C_[3], Sec8_S_[3], Sec8_C_[3] );
HalfAdder sec8ha4( Fir8_S_[5], Fir8_C_[4], Sec8_S_[4], Sec8_C_[4] );
HalfAdder sec8ha5( Fir8_S_[6], Fir8_C_[5], Sec8_S_[5], Sec8_C_[5] );
HalfAdder sec8ha6( Fir8_S_[7], Fir8_C_[6], Sec8_S_[6], Sec8_C_[6] );
HalfAdder sec8ha7( Fir8_S_[8], Fir8_C_[7], Sec8_S_[7], Sec8_C_[7] );
HalfAdder sec8ha8( Fir8_S_[9], Fir8_C_[8], Sec8_S_[8], Sec8_C_[8] );
HalfAdder sec8ha9( Fir8_S_[10], Fir8_C_[9], Sec8_S_[9], Sec8_C_[9] );
HalfAdder sec8ha10( Fir8_S_[11], Fir8_C_[10], Sec8_S_[10], Sec8_C_[10] );
HalfAdder sec8ha11( Fir8_S_[12], Fir8_C_[11], Sec8_S_[11], Sec8_C_[11] );
HalfAdder sec8ha12( Fir8_S_[13], Fir8_C_[12], Sec8_S_[12], Sec8_C_[12] );
HalfAdder sec8ha13( Fir8_S_[14], Fir8_C_[13], Sec8_S_[13], Sec8_C_[13] );
HalfAdder sec8ha14( Fir8_S_[15], Fir8_C_[14], Sec8_S_[14], Sec8_C_[14] );
HalfAdder sec8ha15( Fir8_S_[16], Fir8_C_[15], Sec8_S_[15], Sec8_C_[15] );
HalfAdder sec8ha16( Fir8_S_[17], Fir8_C_[16], Sec8_S_[16], Sec8_C_[16] );
HalfAdder sec8ha17( Fir8_S_[18], Fir8_C_[17], Sec8_S_[17], Sec8_C_[17] );
HalfAdder sec8ha18( Fir8_S_[19], Fir8_C_[18], Sec8_S_[18], Sec8_C_[18] );
HalfAdder sec8ha19( Fir8_S_[20], Fir8_C_[19], Sec8_S_[19], Sec8_C_[19] );
HalfAdder sec8ha20( Fir8_S_[21], Fir8_C_[20], Sec8_S_[20], Sec8_C_[20] );
HalfAdder sec8ha21( Fir8_S_[22], Fir8_C_[21], Sec8_S_[21], Sec8_C_[21] );
HalfAdder sec8ha22( Fir8_S_[23], Fir8_C_[22], Sec8_S_[22], Sec8_C_[22] );
HalfAdder sec8ha23( Fir8_S_[24], Fir8_C_[23], Sec8_S_[23], Sec8_C_[23] );
HalfAdder sec8ha24( Fir8_S_[25], Fir8_C_[24], Sec8_S_[24], Sec8_C_[24] );
HalfAdder sec8ha25( Fir8_S_[26], Fir8_C_[25], Sec8_S_[25], Sec8_C_[25] );
HalfAdder sec8ha26( Fir8_S_[27], Fir8_C_[26], Sec8_S_[26], Sec8_C_[26] );
HalfAdder sec8ha27( Fir8_S_[28], Fir8_C_[27], Sec8_S_[27], Sec8_C_[27] );
HalfAdder sec8ha28( Fir8_S_[29], Fir8_C_[28], Sec8_S_[28], Sec8_C_[28] );
HalfAdder sec8ha29( Fir8_S_[30], Fir8_C_[29], Sec8_S_[29], Sec8_C_[29] );
HalfAdder sec8ha30( Fir8_S_[31], Fir8_C_[30], Sec8_S_[30], Sec8_C_[30] );
HalfAdder sec8ha31( pp23[31], Fir8_C_[31], Sec8_S_[31], Sec8_C_[31] );


HalfAdder sec9ha0( Fir9_S_[1], Fir9_C_[0], Sec9_S_[0], Sec9_C_[0] );
HalfAdder sec9ha1( Fir9_S_[2], Fir9_C_[1], Sec9_S_[1], Sec9_C_[1] );
HalfAdder sec9ha2( Fir9_S_[3], Fir9_C_[2], Sec9_S_[2], Sec9_C_[2] );
HalfAdder sec9ha3( Fir9_S_[4], Fir9_C_[3], Sec9_S_[3], Sec9_C_[3] );
HalfAdder sec9ha4( Fir9_S_[5], Fir9_C_[4], Sec9_S_[4], Sec9_C_[4] );
HalfAdder sec9ha5( Fir9_S_[6], Fir9_C_[5], Sec9_S_[5], Sec9_C_[5] );
HalfAdder sec9ha6( Fir9_S_[7], Fir9_C_[6], Sec9_S_[6], Sec9_C_[6] );
HalfAdder sec9ha7( Fir9_S_[8], Fir9_C_[7], Sec9_S_[7], Sec9_C_[7] );
HalfAdder sec9ha8( Fir9_S_[9], Fir9_C_[8], Sec9_S_[8], Sec9_C_[8] );
HalfAdder sec9ha9( Fir9_S_[10], Fir9_C_[9], Sec9_S_[9], Sec9_C_[9] );
HalfAdder sec9ha10( Fir9_S_[11], Fir9_C_[10], Sec9_S_[10], Sec9_C_[10] );
HalfAdder sec9ha11( Fir9_S_[12], Fir9_C_[11], Sec9_S_[11], Sec9_C_[11] );
HalfAdder sec9ha12( Fir9_S_[13], Fir9_C_[12], Sec9_S_[12], Sec9_C_[12] );
HalfAdder sec9ha13( Fir9_S_[14], Fir9_C_[13], Sec9_S_[13], Sec9_C_[13] );
HalfAdder sec9ha14( Fir9_S_[15], Fir9_C_[14], Sec9_S_[14], Sec9_C_[14] );
HalfAdder sec9ha15( Fir9_S_[16], Fir9_C_[15], Sec9_S_[15], Sec9_C_[15] );
HalfAdder sec9ha16( Fir9_S_[17], Fir9_C_[16], Sec9_S_[16], Sec9_C_[16] );
HalfAdder sec9ha17( Fir9_S_[18], Fir9_C_[17], Sec9_S_[17], Sec9_C_[17] );
HalfAdder sec9ha18( Fir9_S_[19], Fir9_C_[18], Sec9_S_[18], Sec9_C_[18] );
HalfAdder sec9ha19( Fir9_S_[20], Fir9_C_[19], Sec9_S_[19], Sec9_C_[19] );
HalfAdder sec9ha20( Fir9_S_[21], Fir9_C_[20], Sec9_S_[20], Sec9_C_[20] );
HalfAdder sec9ha21( Fir9_S_[22], Fir9_C_[21], Sec9_S_[21], Sec9_C_[21] );
HalfAdder sec9ha22( Fir9_S_[23], Fir9_C_[22], Sec9_S_[22], Sec9_C_[22] );
HalfAdder sec9ha23( Fir9_S_[24], Fir9_C_[23], Sec9_S_[23], Sec9_C_[23] );
HalfAdder sec9ha24( Fir9_S_[25], Fir9_C_[24], Sec9_S_[24], Sec9_C_[24] );
HalfAdder sec9ha25( Fir9_S_[26], Fir9_C_[25], Sec9_S_[25], Sec9_C_[25] );
HalfAdder sec9ha26( Fir9_S_[27], Fir9_C_[26], Sec9_S_[26], Sec9_C_[26] );
HalfAdder sec9ha27( Fir9_S_[28], Fir9_C_[27], Sec9_S_[27], Sec9_C_[27] );
HalfAdder sec9ha28( Fir9_S_[29], Fir9_C_[28], Sec9_S_[28], Sec9_C_[28] );
HalfAdder sec9ha29( Fir9_S_[30], Fir9_C_[29], Sec9_S_[29], Sec9_C_[29] );
HalfAdder sec9ha30( Fir9_S_[31], Fir9_C_[30], Sec9_S_[30], Sec9_C_[30] );
HalfAdder sec9ha31( pp26[31], Fir9_C_[31], Sec9_S_[31], Sec9_C_[31] );

HalfAdder sec10ha0( Fir10_S_[1], Fir10_C_[0], Sec10_S_[0], Sec10_C_[0] );
HalfAdder sec10ha1( Fir10_S_[2], Fir10_C_[1], Sec10_S_[1], Sec10_C_[1] );
HalfAdder sec10ha2( Fir10_S_[3], Fir10_C_[2], Sec10_S_[2], Sec10_C_[2] );
HalfAdder sec10ha3( Fir10_S_[4], Fir10_C_[3], Sec10_S_[3], Sec10_C_[3] );
HalfAdder sec10ha4( Fir10_S_[5], Fir10_C_[4], Sec10_S_[4], Sec10_C_[4] );
HalfAdder sec10ha5( Fir10_S_[6], Fir10_C_[5], Sec10_S_[5], Sec10_C_[5] );
HalfAdder sec10ha6( Fir10_S_[7], Fir10_C_[6], Sec10_S_[6], Sec10_C_[6] );
HalfAdder sec10ha7( Fir10_S_[8], Fir10_C_[7], Sec10_S_[7], Sec10_C_[7] );
HalfAdder sec10ha8( Fir10_S_[9], Fir10_C_[8], Sec10_S_[8], Sec10_C_[8] );
HalfAdder sec10ha9( Fir10_S_[10], Fir10_C_[9], Sec10_S_[9], Sec10_C_[9] );
HalfAdder sec10ha10( Fir10_S_[11], Fir10_C_[10], Sec10_S_[10], Sec10_C_[10] );
HalfAdder sec10ha11( Fir10_S_[12], Fir10_C_[11], Sec10_S_[11], Sec10_C_[11] );
HalfAdder sec10ha12( Fir10_S_[13], Fir10_C_[12], Sec10_S_[12], Sec10_C_[12] );
HalfAdder sec10ha13( Fir10_S_[14], Fir10_C_[13], Sec10_S_[13], Sec10_C_[13] );
HalfAdder sec10ha14( Fir10_S_[15], Fir10_C_[14], Sec10_S_[14], Sec10_C_[14] );
HalfAdder sec10ha15( Fir10_S_[16], Fir10_C_[15], Sec10_S_[15], Sec10_C_[15] );
HalfAdder sec10ha16( Fir10_S_[17], Fir10_C_[16], Sec10_S_[16], Sec10_C_[16] );
HalfAdder sec10ha17( Fir10_S_[18], Fir10_C_[17], Sec10_S_[17], Sec10_C_[17] );
HalfAdder sec10ha18( Fir10_S_[19], Fir10_C_[18], Sec10_S_[18], Sec10_C_[18] );
HalfAdder sec10ha19( Fir10_S_[20], Fir10_C_[19], Sec10_S_[19], Sec10_C_[19] );
HalfAdder sec10ha20( Fir10_S_[21], Fir10_C_[20], Sec10_S_[20], Sec10_C_[20] );
HalfAdder sec10ha21( Fir10_S_[22], Fir10_C_[21], Sec10_S_[21], Sec10_C_[21] );
HalfAdder sec10ha22( Fir10_S_[23], Fir10_C_[22], Sec10_S_[22], Sec10_C_[22] );
HalfAdder sec10ha23( Fir10_S_[24], Fir10_C_[23], Sec10_S_[23], Sec10_C_[23] );
HalfAdder sec10ha24( Fir10_S_[25], Fir10_C_[24], Sec10_S_[24], Sec10_C_[24] );
HalfAdder sec10ha25( Fir10_S_[26], Fir10_C_[25], Sec10_S_[25], Sec10_C_[25] );
HalfAdder sec10ha26( Fir10_S_[27], Fir10_C_[26], Sec10_S_[26], Sec10_C_[26] );
HalfAdder sec10ha27( Fir10_S_[28], Fir10_C_[27], Sec10_S_[27], Sec10_C_[27] );
HalfAdder sec10ha28( Fir10_S_[29], Fir10_C_[28], Sec10_S_[28], Sec10_C_[28] );
HalfAdder sec10ha29( Fir10_S_[30], Fir10_C_[29], Sec10_S_[29], Sec10_C_[29] );
HalfAdder sec10ha30( Fir10_S_[31], Fir10_C_[30], Sec10_S_[30], Sec10_C_[30] );
HalfAdder sec10ha31( pp29[31], Fir10_C_[31], Sec10_S_[31], Sec10_C_[31] );


HalfAdder sec11ha0( Fir11_S_[1], Fir11_C_[0], Sec11_S_[0], Sec11_C_[0] );
HalfAdder sec11ha1( Fir11_S_[2], Fir11_C_[1], Sec11_S_[1], Sec11_C_[1] );
HalfAdder sec11ha2( Fir11_S_[3], Fir11_C_[2], Sec11_S_[2], Sec11_C_[2] );
HalfAdder sec11ha3( Fir11_S_[4], Fir11_C_[3], Sec11_S_[3], Sec11_C_[3] );
HalfAdder sec11ha4( Fir11_S_[5], Fir11_C_[4], Sec11_S_[4], Sec11_C_[4] );
HalfAdder sec11ha5( Fir11_S_[6], Fir11_C_[5], Sec11_S_[5], Sec11_C_[5] );
HalfAdder sec11ha6( Fir11_S_[7], Fir11_C_[6], Sec11_S_[6], Sec11_C_[6] );
HalfAdder sec11ha7( Fir11_S_[8], Fir11_C_[7], Sec11_S_[7], Sec11_C_[7] );
HalfAdder sec11ha8( Fir11_S_[9], Fir11_C_[8], Sec11_S_[8], Sec11_C_[8] );
HalfAdder sec11ha9( Fir11_S_[10], Fir11_C_[9], Sec11_S_[9], Sec11_C_[9] );
HalfAdder sec11ha10( Fir11_S_[11], Fir11_C_[10], Sec11_S_[10], Sec11_C_[10] );
HalfAdder sec11ha11( Fir11_S_[12], Fir11_C_[11], Sec11_S_[11], Sec11_C_[11] );
HalfAdder sec11ha12( Fir11_S_[13], Fir11_C_[12], Sec11_S_[12], Sec11_C_[12] );
HalfAdder sec11ha13( Fir11_S_[14], Fir11_C_[13], Sec11_S_[13], Sec11_C_[13] );
HalfAdder sec11ha14( Fir11_S_[15], Fir11_C_[14], Sec11_S_[14], Sec11_C_[14] );
HalfAdder sec11ha15( Fir11_S_[16], Fir11_C_[15], Sec11_S_[15], Sec11_C_[15] );
HalfAdder sec11ha16( Fir11_S_[17], Fir11_C_[16], Sec11_S_[16], Sec11_C_[16] );
HalfAdder sec11ha17( Fir11_S_[18], Fir11_C_[17], Sec11_S_[17], Sec11_C_[17] );
HalfAdder sec11ha18( Fir11_S_[19], Fir11_C_[18], Sec11_S_[18], Sec11_C_[18] );
HalfAdder sec11ha19( Fir11_S_[20], Fir11_C_[19], Sec11_S_[19], Sec11_C_[19] );
HalfAdder sec11ha20( Fir11_S_[21], Fir11_C_[20], Sec11_S_[20], Sec11_C_[20] );
HalfAdder sec11ha21( Fir11_S_[22], Fir11_C_[21], Sec11_S_[21], Sec11_C_[21] );
HalfAdder sec11ha22( Fir11_S_[23], Fir11_C_[22], Sec11_S_[22], Sec11_C_[22] );
HalfAdder sec11ha23( Fir11_S_[24], Fir11_C_[23], Sec11_S_[23], Sec11_C_[23] );
HalfAdder sec11ha24( Fir11_S_[25], Fir11_C_[24], Sec11_S_[24], Sec11_C_[24] );
HalfAdder sec11ha25( Fir11_S_[26], Fir11_C_[25], Sec11_S_[25], Sec11_C_[25] );
HalfAdder sec11ha26( Fir11_S_[27], Fir11_C_[26], Sec11_S_[26], Sec11_C_[26] );
HalfAdder sec11ha27( Fir11_S_[28], Fir11_C_[27], Sec11_S_[27], Sec11_C_[27] );
HalfAdder sec11ha28( Fir11_S_[29], Fir11_C_[28], Sec11_S_[28], Sec11_C_[28] );
HalfAdder sec11ha29( Fir11_S_[30], Fir11_C_[29], Sec11_S_[29], Sec11_C_[29] );
HalfAdder sec11ha30( pp31[31], Fir11_C_[30], Sec11_S_[30], Sec11_C_[30] );



reg	[31: 0]	Sec1_S, Sec1_C;
reg	[31: 0]	Sec2_S, Sec2_C;
reg	[31: 0]	Sec3_S, Sec3_C;
reg	[31: 0]	Sec4_S, Sec4_C;
reg	[31: 0]	Sec5_S, Sec5_C;
reg	[31: 0]	Sec6_S, Sec6_C;
reg	[31: 0]	Sec7_S, Sec7_C;
reg	[31: 0]	Sec8_S, Sec8_C;
reg	[31: 0]	Sec9_S, Sec9_C;
reg	[31: 0]	Sec10_S, Sec10_C;
reg	[30: 0]	Sec11_S, Sec11_C;
reg done1;
reg state_done1;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Sec1_S  <= 32'b0;  Sec1_C  <= 32'b0;
        Sec2_S  <= 32'b0;  Sec2_C  <= 32'b0;
        Sec3_S  <= 32'b0;  Sec3_C  <= 32'b0;
        Sec4_S  <= 32'b0;  Sec4_C  <= 32'b0;
        Sec5_S  <= 32'b0;  Sec5_C  <= 32'b0;
        Sec6_S  <= 32'b0;  Sec6_C  <= 32'b0;
        Sec7_S  <= 32'b0;  Sec7_C  <= 32'b0;
        Sec8_S  <= 32'b0;  Sec8_C  <= 32'b0;
        Sec9_S  <= 32'b0;  Sec9_C  <= 32'b0;
        Sec10_S <= 32'b0;  Sec10_C <= 32'b0;
        Sec11_S <= 31'b0;  Sec11_C <= 31'b0;
        done1       <= 1'b0;
        state_done1 <= 1'b0;
    end
    else begin
        case (state_done1)
            1'b0: begin
                if (done0) begin
                    Sec1_S  <= Sec1_S_; Sec1_C  <= Sec1_C_;
                    Sec2_S  <= Sec2_S_; Sec2_C  <= Sec2_C_;
                    Sec3_S  <= Sec3_S_; Sec3_C  <= Sec3_C_;
                    Sec4_S  <= Sec4_S_; Sec4_C  <= Sec4_C_;
                    Sec5_S  <= Sec5_S_; Sec5_C  <= Sec5_C_;
                    Sec6_S  <= Sec6_S_; Sec6_C  <= Sec6_C_;
                    Sec7_S  <= Sec7_S_; Sec7_C  <= Sec7_C_;
                    Sec8_S  <= Sec8_S_; Sec8_C  <= Sec8_C_;
                    Sec9_S  <= Sec9_S_; Sec9_C  <= Sec9_C_;
                    Sec10_S <= Sec10_S_; Sec10_C <= Sec10_C_;
                    Sec11_S <= Sec11_S_; Sec11_C <= Sec11_C_;
                    done1 <= 1'b1;
                    state_done1 <= 1'b1;
                end else begin
                    done1 <= 1'b0;
                end
            end
            1'b1: begin
                done1 <= 1'b0;
                if (!done0)
                    state_done1 <= 1'b0;
            end
        endcase
    end
end
//===================Third stage===============================

wire	[31: 0]	Thi1_S, Thi1_C;
wire	[33: 0]	Thi2_S, Thi2_C;
wire	[31: 0]	Thi3_S, Thi3_C;
wire	[33: 0]	Thi4_S, Thi4_C;
wire	[31: 0]	Thi5_S, Thi5_C;
wire	[33: 0]	Thi6_S, Thi6_C;
wire	[31: 0]	Thi7_S, Thi7_C;


FullAdder thi1fa1( Sec1_C[0], Sec1_S[1], pp3[0], Thi1_S[0], Thi1_C[0] );
FullAdder thi1fa2( Sec1_C[1], Sec1_S[2], Fir2_S_[0], Thi1_S[1], Thi1_C[1] );
FullAdder thi1fa3( Sec1_C[2], Sec1_S[3], Sec2_S[0], Thi1_S[2], Thi1_C[2] );
FullAdder thi1fa4( Sec1_C[3], Sec1_S[4], Sec2_S[1], Thi1_S[3], Thi1_C[3] );
FullAdder thi1fa5( Sec1_C[4], Sec1_S[5], Sec2_S[2], Thi1_S[4], Thi1_C[4] );
FullAdder thi1fa6( Sec1_C[5], Sec1_S[6], Sec2_S[3], Thi1_S[5], Thi1_C[5] );
FullAdder thi1fa7( Sec1_C[6], Sec1_S[7], Sec2_S[4], Thi1_S[6], Thi1_C[6] );
FullAdder thi1fa8( Sec1_C[7], Sec1_S[8], Sec2_S[5], Thi1_S[7], Thi1_C[7] );
FullAdder thi1fa9( Sec1_C[8], Sec1_S[9], Sec2_S[6], Thi1_S[8], Thi1_C[8] );
FullAdder thi1fa10( Sec1_C[9], Sec1_S[10], Sec2_S[7], Thi1_S[9], Thi1_C[9] );
FullAdder thi1fa11( Sec1_C[10], Sec1_S[11], Sec2_S[8], Thi1_S[10], Thi1_C[10] );
FullAdder thi1fa12( Sec1_C[11], Sec1_S[12], Sec2_S[9], Thi1_S[11], Thi1_C[11] );
FullAdder thi1fa13( Sec1_C[12], Sec1_S[13], Sec2_S[10], Thi1_S[12], Thi1_C[12] );
FullAdder thi1fa14( Sec1_C[13], Sec1_S[14], Sec2_S[11], Thi1_S[13], Thi1_C[13] );
FullAdder thi1fa15( Sec1_C[14], Sec1_S[15], Sec2_S[12], Thi1_S[14], Thi1_C[14] );
FullAdder thi1fa16( Sec1_C[15], Sec1_S[16], Sec2_S[13], Thi1_S[15], Thi1_C[15] );
FullAdder thi1fa17( Sec1_C[16], Sec1_S[17], Sec2_S[14], Thi1_S[16], Thi1_C[16] );
FullAdder thi1fa18( Sec1_C[17], Sec1_S[18], Sec2_S[15], Thi1_S[17], Thi1_C[17] );
FullAdder thi1fa19( Sec1_C[18], Sec1_S[19], Sec2_S[16], Thi1_S[18], Thi1_C[18] );
FullAdder thi1fa20( Sec1_C[19], Sec1_S[20], Sec2_S[17], Thi1_S[19], Thi1_C[19] );
FullAdder thi1fa21( Sec1_C[20], Sec1_S[21], Sec2_S[18], Thi1_S[20], Thi1_C[20] );
FullAdder thi1fa22( Sec1_C[21], Sec1_S[22], Sec2_S[19], Thi1_S[21], Thi1_C[21] );
FullAdder thi1fa23( Sec1_C[22], Sec1_S[23], Sec2_S[20], Thi1_S[22], Thi1_C[22] );
FullAdder thi1fa24( Sec1_C[23], Sec1_S[24], Sec2_S[21], Thi1_S[23], Thi1_C[23] );
FullAdder thi1fa25( Sec1_C[24], Sec1_S[25], Sec2_S[22], Thi1_S[24], Thi1_C[24] );
FullAdder thi1fa26( Sec1_C[25], Sec1_S[26], Sec2_S[23], Thi1_S[25], Thi1_C[25] );
FullAdder thi1fa27( Sec1_C[26], Sec1_S[27], Sec2_S[24], Thi1_S[26], Thi1_C[26] );
FullAdder thi1fa28( Sec1_C[27], Sec1_S[28], Sec2_S[25], Thi1_S[27], Thi1_C[27] );
FullAdder thi1fa29( Sec1_C[28], Sec1_S[29], Sec2_S[26], Thi1_S[28], Thi1_C[28] );
FullAdder thi1fa30( Sec1_C[29], Sec1_S[30], Sec2_S[27], Thi1_S[29], Thi1_C[29] );
FullAdder thi1fa31( Sec1_C[30], Sec1_S[31], Sec2_S[28], Thi1_S[30], Thi1_C[30] );
HalfAdder thi1fa32( Sec1_C[31], Sec2_S[29], Thi1_S[31], Thi1_C[31] );


HalfAdder thi2fa1( Sec2_C[0], pp6[0], Thi2_S[0], Thi2_C[0] );
HalfAdder thi2fa2( Sec2_C[1], Fir3_S_[0], Thi2_S[1], Thi2_C[1] );
HalfAdder thi2fa3( Sec2_C[2], Sec3_S[0], Thi2_S[2], Thi2_C[2] );
FullAdder thi2fa4( Sec2_C[3], Sec3_S[1], Sec3_C[0], Thi2_S[3], Thi2_C[3] );
FullAdder thi2fa5( Sec2_C[4], Sec3_S[2], Sec3_C[1], Thi2_S[4], Thi2_C[4] );
FullAdder thi2fa6( Sec2_C[5], Sec3_S[3], Sec3_C[2], Thi2_S[5], Thi2_C[5] );
FullAdder thi2fa7( Sec2_C[6], Sec3_S[4], Sec3_C[3], Thi2_S[6], Thi2_C[6] );
FullAdder thi2fa8( Sec2_C[7], Sec3_S[5], Sec3_C[4], Thi2_S[7], Thi2_C[7] );
FullAdder thi2fa9( Sec2_C[8], Sec3_S[6], Sec3_C[5], Thi2_S[8], Thi2_C[8] );
FullAdder thi2fa10( Sec2_C[9], Sec3_S[7], Sec3_C[6], Thi2_S[9], Thi2_C[9] );
FullAdder thi2fa11( Sec2_C[10], Sec3_S[8], Sec3_C[7], Thi2_S[10], Thi2_C[10] );
FullAdder thi2fa12( Sec2_C[11], Sec3_S[9], Sec3_C[8], Thi2_S[11], Thi2_C[11] );
FullAdder thi2fa13( Sec2_C[12], Sec3_S[10], Sec3_C[9], Thi2_S[12], Thi2_C[12] );
FullAdder thi2fa14( Sec2_C[13], Sec3_S[11], Sec3_C[10], Thi2_S[13], Thi2_C[13] );
FullAdder thi2fa15( Sec2_C[14], Sec3_S[12], Sec3_C[11], Thi2_S[14], Thi2_C[14] );
FullAdder thi2fa16( Sec2_C[15], Sec3_S[13], Sec3_C[12], Thi2_S[15], Thi2_C[15] );
FullAdder thi2fa17( Sec2_C[16], Sec3_S[14], Sec3_C[13], Thi2_S[16], Thi2_C[16] );
FullAdder thi2fa18( Sec2_C[17], Sec3_S[15], Sec3_C[14], Thi2_S[17], Thi2_C[17] );
FullAdder thi2fa19( Sec2_C[18], Sec3_S[16], Sec3_C[15], Thi2_S[18], Thi2_C[18] );
FullAdder thi2fa20( Sec2_C[19], Sec3_S[17], Sec3_C[16], Thi2_S[19], Thi2_C[19] );
FullAdder thi2fa21( Sec2_C[20], Sec3_S[18], Sec3_C[17], Thi2_S[20], Thi2_C[20] );
FullAdder thi2fa22( Sec2_C[21], Sec3_S[19], Sec3_C[18], Thi2_S[21], Thi2_C[21] );
FullAdder thi2fa23( Sec2_C[22], Sec3_S[20], Sec3_C[19], Thi2_S[22], Thi2_C[22] );
FullAdder thi2fa24( Sec2_C[23], Sec3_S[21], Sec3_C[20], Thi2_S[23], Thi2_C[23] );
FullAdder thi2fa25( Sec2_C[24], Sec3_S[22], Sec3_C[21], Thi2_S[24], Thi2_C[24] );
FullAdder thi2fa26( Sec2_C[25], Sec3_S[23], Sec3_C[22], Thi2_S[25], Thi2_C[25] );
FullAdder thi2fa27( Sec2_C[26], Sec3_S[24], Sec3_C[23], Thi2_S[26], Thi2_C[26] );
FullAdder thi2fa28( Sec2_C[27], Sec3_S[25], Sec3_C[24], Thi2_S[27], Thi2_C[27] );
FullAdder thi2fa29( Sec2_C[28], Sec3_S[26], Sec3_C[25], Thi2_S[28], Thi2_C[28] );
FullAdder thi2fa30( Sec2_C[29], Sec3_S[27], Sec3_C[26], Thi2_S[29], Thi2_C[29] );
FullAdder thi2fa31( Sec2_C[30], Sec3_S[28], Sec3_C[27], Thi2_S[30], Thi2_C[30] );
FullAdder thi2fa32( Sec2_C[31], Sec3_S[29], Sec3_C[28], Thi2_S[31], Thi2_C[31] );
HalfAdder thi2fa33( Sec3_S[30], Sec3_C[29], Thi2_S[32], Thi2_C[32]);
HalfAdder thi2fa34( Sec3_S[31], Sec3_C[30], Thi2_S[33], Thi2_C[33]);

FullAdder thi3fa1( Sec4_C[0], Sec4_S[1], pp12[0], Thi3_S[0], Thi3_C[0] );
FullAdder thi3fa2( Sec4_C[1], Sec4_S[2], Fir5_S_[0], Thi3_S[1], Thi3_C[1] );
FullAdder thi3fa3( Sec4_C[2], Sec4_S[3], Sec5_S[0], Thi3_S[2], Thi3_C[2] );
FullAdder thi3fa4( Sec4_C[3], Sec4_S[4], Sec5_S[1], Thi3_S[3], Thi3_C[3] );
FullAdder thi3fa5( Sec4_C[4], Sec4_S[5], Sec5_S[2], Thi3_S[4], Thi3_C[4] );
FullAdder thi3fa6( Sec4_C[5], Sec4_S[6], Sec5_S[3], Thi3_S[5], Thi3_C[5] );
FullAdder thi3fa7( Sec4_C[6], Sec4_S[7], Sec5_S[4], Thi3_S[6], Thi3_C[6] );
FullAdder thi3fa8( Sec4_C[7], Sec4_S[8], Sec5_S[5], Thi3_S[7], Thi3_C[7] );
FullAdder thi3fa9( Sec4_C[8], Sec4_S[9], Sec5_S[6], Thi3_S[8], Thi3_C[8] );
FullAdder thi3fa10( Sec4_C[9], Sec4_S[10], Sec5_S[7], Thi3_S[9], Thi3_C[9] );
FullAdder thi3fa11( Sec4_C[10], Sec4_S[11], Sec5_S[8], Thi3_S[10], Thi3_C[10] );
FullAdder thi3fa12( Sec4_C[11], Sec4_S[12], Sec5_S[9], Thi3_S[11], Thi3_C[11] );
FullAdder thi3fa13( Sec4_C[12], Sec4_S[13], Sec5_S[10], Thi3_S[12], Thi3_C[12] );
FullAdder thi3fa14( Sec4_C[13], Sec4_S[14], Sec5_S[11], Thi3_S[13], Thi3_C[13] );
FullAdder thi3fa15( Sec4_C[14], Sec4_S[15], Sec5_S[12], Thi3_S[14], Thi3_C[14] );
FullAdder thi3fa16( Sec4_C[15], Sec4_S[16], Sec5_S[13], Thi3_S[15], Thi3_C[15] );
FullAdder thi3fa17( Sec4_C[16], Sec4_S[17], Sec5_S[14], Thi3_S[16], Thi3_C[16] );
FullAdder thi3fa18( Sec4_C[17], Sec4_S[18], Sec5_S[15], Thi3_S[17], Thi3_C[17] );
FullAdder thi3fa19( Sec4_C[18], Sec4_S[19], Sec5_S[16], Thi3_S[18], Thi3_C[18] );
FullAdder thi3fa20( Sec4_C[19], Sec4_S[20], Sec5_S[17], Thi3_S[19], Thi3_C[19] );
FullAdder thi3fa21( Sec4_C[20], Sec4_S[21], Sec5_S[18], Thi3_S[20], Thi3_C[20] );
FullAdder thi3fa22( Sec4_C[21], Sec4_S[22], Sec5_S[19], Thi3_S[21], Thi3_C[21] );
FullAdder thi3fa23( Sec4_C[22], Sec4_S[23], Sec5_S[20], Thi3_S[22], Thi3_C[22] );
FullAdder thi3fa24( Sec4_C[23], Sec4_S[24], Sec5_S[21], Thi3_S[23], Thi3_C[23] );
FullAdder thi3fa25( Sec4_C[24], Sec4_S[25], Sec5_S[22], Thi3_S[24], Thi3_C[24] );
FullAdder thi3fa26( Sec4_C[25], Sec4_S[26], Sec5_S[23], Thi3_S[25], Thi3_C[25] );
FullAdder thi3fa27( Sec4_C[26], Sec4_S[27], Sec5_S[24], Thi3_S[26], Thi3_C[26] );
FullAdder thi3fa28( Sec4_C[27], Sec4_S[28], Sec5_S[25], Thi3_S[27], Thi3_C[27] );
FullAdder thi3fa29( Sec4_C[28], Sec4_S[29], Sec5_S[26], Thi3_S[28], Thi3_C[28] );
FullAdder thi3fa30( Sec4_C[29], Sec4_S[30], Sec5_S[27], Thi3_S[29], Thi3_C[29] );
FullAdder thi3fa31( Sec4_C[30], Sec4_S[31], Sec5_S[28], Thi3_S[30], Thi3_C[30] );
HalfAdder thi3fa32( Sec4_C[31], Sec5_S[29], Thi3_S[31], Thi3_C[31] );


HalfAdder thi4fa1( Sec5_C[0], pp15[0], Thi4_S[0], Thi4_C[0] );
HalfAdder thi4fa2( Sec5_C[1], Fir6_S_[0], Thi4_S[1], Thi4_C[1] );
HalfAdder thi4fa3( Sec5_C[2], Sec6_S[0], Thi4_S[2], Thi4_C[2] );
FullAdder thi4fa4( Sec5_C[3], Sec6_S[1], Sec6_C[0], Thi4_S[3], Thi4_C[3] );
FullAdder thi4fa5( Sec5_C[4], Sec6_S[2], Sec6_C[1], Thi4_S[4], Thi4_C[4] );
FullAdder thi4fa6( Sec5_C[5], Sec6_S[3], Sec6_C[2], Thi4_S[5], Thi4_C[5] );
FullAdder thi4fa7( Sec5_C[6], Sec6_S[4], Sec6_C[3], Thi4_S[6], Thi4_C[6] );
FullAdder thi4fa8( Sec5_C[7], Sec6_S[5], Sec6_C[4], Thi4_S[7], Thi4_C[7] );
FullAdder thi4fa9( Sec5_C[8], Sec6_S[6], Sec6_C[5], Thi4_S[8], Thi4_C[8] );
FullAdder thi4fa10( Sec5_C[9], Sec6_S[7], Sec6_C[6], Thi4_S[9], Thi4_C[9] );
FullAdder thi4fa11( Sec5_C[10], Sec6_S[8], Sec6_C[7], Thi4_S[10], Thi4_C[10] );
FullAdder thi4fa12( Sec5_C[11], Sec6_S[9], Sec6_C[8], Thi4_S[11], Thi4_C[11] );
FullAdder thi4fa13( Sec5_C[12], Sec6_S[10], Sec6_C[9], Thi4_S[12], Thi4_C[12] );
FullAdder thi4fa14( Sec5_C[13], Sec6_S[11], Sec6_C[10], Thi4_S[13], Thi4_C[13] );
FullAdder thi4fa15( Sec5_C[14], Sec6_S[12], Sec6_C[11], Thi4_S[14], Thi4_C[14] );
FullAdder thi4fa16( Sec5_C[15], Sec6_S[13], Sec6_C[12], Thi4_S[15], Thi4_C[15] );
FullAdder thi4fa17( Sec5_C[16], Sec6_S[14], Sec6_C[13], Thi4_S[16], Thi4_C[16] );
FullAdder thi4fa18( Sec5_C[17], Sec6_S[15], Sec6_C[14], Thi4_S[17], Thi4_C[17] );
FullAdder thi4fa19( Sec5_C[18], Sec6_S[16], Sec6_C[15], Thi4_S[18], Thi4_C[18] );
FullAdder thi4fa20( Sec5_C[19], Sec6_S[17], Sec6_C[16], Thi4_S[19], Thi4_C[19] );
FullAdder thi4fa21( Sec5_C[20], Sec6_S[18], Sec6_C[17], Thi4_S[20], Thi4_C[20] );
FullAdder thi4fa22( Sec5_C[21], Sec6_S[19], Sec6_C[18], Thi4_S[21], Thi4_C[21] );
FullAdder thi4fa23( Sec5_C[22], Sec6_S[20], Sec6_C[19], Thi4_S[22], Thi4_C[22] );
FullAdder thi4fa24( Sec5_C[23], Sec6_S[21], Sec6_C[20], Thi4_S[23], Thi4_C[23] );
FullAdder thi4fa25( Sec5_C[24], Sec6_S[22], Sec6_C[21], Thi4_S[24], Thi4_C[24] );
FullAdder thi4fa26( Sec5_C[25], Sec6_S[23], Sec6_C[22], Thi4_S[25], Thi4_C[25] );
FullAdder thi4fa27( Sec5_C[26], Sec6_S[24], Sec6_C[23], Thi4_S[26], Thi4_C[26] );
FullAdder thi4fa28( Sec5_C[27], Sec6_S[25], Sec6_C[24], Thi4_S[27], Thi4_C[27] );
FullAdder thi4fa29( Sec5_C[28], Sec6_S[26], Sec6_C[25], Thi4_S[28], Thi4_C[28] );
FullAdder thi4fa30( Sec5_C[29], Sec6_S[27], Sec6_C[26], Thi4_S[29], Thi4_C[29] );
FullAdder thi4fa31( Sec5_C[30], Sec6_S[28], Sec6_C[27], Thi4_S[30], Thi4_C[30] );
FullAdder thi4fa32( Sec5_C[31], Sec6_S[29], Sec6_C[28], Thi4_S[31], Thi4_C[31] );
HalfAdder thi4fa33( Sec6_S[30], Sec6_C[29], Thi4_S[32], Thi4_C[32]);
HalfAdder thi4fa34( Sec6_S[31], Sec6_C[30], Thi4_S[33], Thi4_C[33]);

FullAdder thi5fa1( Sec7_C[0], Sec7_S[1], pp21[0], Thi5_S[0], Thi5_C[0] );
FullAdder thi5fa2( Sec7_C[1], Sec7_S[2], Fir8_S_[0], Thi5_S[1], Thi5_C[1] );
FullAdder thi5fa3( Sec7_C[2], Sec7_S[3], Sec8_S[0], Thi5_S[2], Thi5_C[2] );
FullAdder thi5fa4( Sec7_C[3], Sec7_S[4], Sec8_S[1], Thi5_S[3], Thi5_C[3] );
FullAdder thi5fa5( Sec7_C[4], Sec7_S[5], Sec8_S[2], Thi5_S[4], Thi5_C[4] );
FullAdder thi5fa6( Sec7_C[5], Sec7_S[6], Sec8_S[3], Thi5_S[5], Thi5_C[5] );
FullAdder thi5fa7( Sec7_C[6], Sec7_S[7], Sec8_S[4], Thi5_S[6], Thi5_C[6] );
FullAdder thi5fa8( Sec7_C[7], Sec7_S[8], Sec8_S[5], Thi5_S[7], Thi5_C[7] );
FullAdder thi5fa9( Sec7_C[8], Sec7_S[9], Sec8_S[6], Thi5_S[8], Thi5_C[8] );
FullAdder thi5fa10( Sec7_C[9], Sec7_S[10], Sec8_S[7], Thi5_S[9], Thi5_C[9] );
FullAdder thi5fa11( Sec7_C[10], Sec7_S[11], Sec8_S[8], Thi5_S[10], Thi5_C[10] );
FullAdder thi5fa12( Sec7_C[11], Sec7_S[12], Sec8_S[9], Thi5_S[11], Thi5_C[11] );
FullAdder thi5fa13( Sec7_C[12], Sec7_S[13], Sec8_S[10], Thi5_S[12], Thi5_C[12] );
FullAdder thi5fa14( Sec7_C[13], Sec7_S[14], Sec8_S[11], Thi5_S[13], Thi5_C[13] );
FullAdder thi5fa15( Sec7_C[14], Sec7_S[15], Sec8_S[12], Thi5_S[14], Thi5_C[14] );
FullAdder thi5fa16( Sec7_C[15], Sec7_S[16], Sec8_S[13], Thi5_S[15], Thi5_C[15] );
FullAdder thi5fa17( Sec7_C[16], Sec7_S[17], Sec8_S[14], Thi5_S[16], Thi5_C[16] );
FullAdder thi5fa18( Sec7_C[17], Sec7_S[18], Sec8_S[15], Thi5_S[17], Thi5_C[17] );
FullAdder thi5fa19( Sec7_C[18], Sec7_S[19], Sec8_S[16], Thi5_S[18], Thi5_C[18] );
FullAdder thi5fa20( Sec7_C[19], Sec7_S[20], Sec8_S[17], Thi5_S[19], Thi5_C[19] );
FullAdder thi5fa21( Sec7_C[20], Sec7_S[21], Sec8_S[18], Thi5_S[20], Thi5_C[20] );
FullAdder thi5fa22( Sec7_C[21], Sec7_S[22], Sec8_S[19], Thi5_S[21], Thi5_C[21] );
FullAdder thi5fa23( Sec7_C[22], Sec7_S[23], Sec8_S[20], Thi5_S[22], Thi5_C[22] );
FullAdder thi5fa24( Sec7_C[23], Sec7_S[24], Sec8_S[21], Thi5_S[23], Thi5_C[23] );
FullAdder thi5fa25( Sec7_C[24], Sec7_S[25], Sec8_S[22], Thi5_S[24], Thi5_C[24] );
FullAdder thi5fa26( Sec7_C[25], Sec7_S[26], Sec8_S[23], Thi5_S[25], Thi5_C[25] );
FullAdder thi5fa27( Sec7_C[26], Sec7_S[27], Sec8_S[24], Thi5_S[26], Thi5_C[26] );
FullAdder thi5fa28( Sec7_C[27], Sec7_S[28], Sec8_S[25], Thi5_S[27], Thi5_C[27] );
FullAdder thi5fa29( Sec7_C[28], Sec7_S[29], Sec8_S[26], Thi5_S[28], Thi5_C[28] );
FullAdder thi5fa30( Sec7_C[29], Sec7_S[30], Sec8_S[27], Thi5_S[29], Thi5_C[29] );
FullAdder thi5fa31( Sec7_C[30], Sec7_S[31], Sec8_S[28], Thi5_S[30], Thi5_C[30] );
HalfAdder thi5fa32( Sec7_C[31], Sec8_S[29], Thi5_S[31], Thi5_C[31] );

HalfAdder thi6fa1( Sec8_C[0], pp24[0], Thi6_S[0], Thi6_C[0] );
HalfAdder thi6fa2( Sec8_C[1], Fir9_S_[0], Thi6_S[1], Thi6_C[1] );
HalfAdder thi6fa3( Sec8_C[2], Sec9_S[0], Thi6_S[2], Thi6_C[2] );
FullAdder thi6fa4( Sec8_C[3], Sec9_S[1], Sec9_C[0], Thi6_S[3], Thi6_C[3] );
FullAdder thi6fa5( Sec8_C[4], Sec9_S[2], Sec9_C[1], Thi6_S[4], Thi6_C[4] );
FullAdder thi6fa6( Sec8_C[5], Sec9_S[3], Sec9_C[2], Thi6_S[5], Thi6_C[5] );
FullAdder thi6fa7( Sec8_C[6], Sec9_S[4], Sec9_C[3], Thi6_S[6], Thi6_C[6] );
FullAdder thi6fa8( Sec8_C[7], Sec9_S[5], Sec9_C[4], Thi6_S[7], Thi6_C[7] );
FullAdder thi6fa9( Sec8_C[8], Sec9_S[6], Sec9_C[5], Thi6_S[8], Thi6_C[8] );
FullAdder thi6fa10( Sec8_C[9], Sec9_S[7], Sec9_C[6], Thi6_S[9], Thi6_C[9] );
FullAdder thi6fa11( Sec8_C[10], Sec9_S[8], Sec9_C[7], Thi6_S[10], Thi6_C[10] );
FullAdder thi6fa12( Sec8_C[11], Sec9_S[9], Sec9_C[8], Thi6_S[11], Thi6_C[11] );
FullAdder thi6fa13( Sec8_C[12], Sec9_S[10], Sec9_C[9], Thi6_S[12], Thi6_C[12] );
FullAdder thi6fa14( Sec8_C[13], Sec9_S[11], Sec9_C[10], Thi6_S[13], Thi6_C[13] );
FullAdder thi6fa15( Sec8_C[14], Sec9_S[12], Sec9_C[11], Thi6_S[14], Thi6_C[14] );
FullAdder thi6fa16( Sec8_C[15], Sec9_S[13], Sec9_C[12], Thi6_S[15], Thi6_C[15] );
FullAdder thi6fa17( Sec8_C[16], Sec9_S[14], Sec9_C[13], Thi6_S[16], Thi6_C[16] );
FullAdder thi6fa18( Sec8_C[17], Sec9_S[15], Sec9_C[14], Thi6_S[17], Thi6_C[17] );
FullAdder thi6fa19( Sec8_C[18], Sec9_S[16], Sec9_C[15], Thi6_S[18], Thi6_C[18] );
FullAdder thi6fa20( Sec8_C[19], Sec9_S[17], Sec9_C[16], Thi6_S[19], Thi6_C[19] );
FullAdder thi6fa21( Sec8_C[20], Sec9_S[18], Sec9_C[17], Thi6_S[20], Thi6_C[20] );
FullAdder thi6fa22( Sec8_C[21], Sec9_S[19], Sec9_C[18], Thi6_S[21], Thi6_C[21] );
FullAdder thi6fa23( Sec8_C[22], Sec9_S[20], Sec9_C[19], Thi6_S[22], Thi6_C[22] );
FullAdder thi6fa24( Sec8_C[23], Sec9_S[21], Sec9_C[20], Thi6_S[23], Thi6_C[23] );
FullAdder thi6fa25( Sec8_C[24], Sec9_S[22], Sec9_C[21], Thi6_S[24], Thi6_C[24] );
FullAdder thi6fa26( Sec8_C[25], Sec9_S[23], Sec9_C[22], Thi6_S[25], Thi6_C[25] );
FullAdder thi6fa27( Sec8_C[26], Sec9_S[24], Sec9_C[23], Thi6_S[26], Thi6_C[26] );
FullAdder thi6fa28( Sec8_C[27], Sec9_S[25], Sec9_C[24], Thi6_S[27], Thi6_C[27] );
FullAdder thi6fa29( Sec8_C[28], Sec9_S[26], Sec9_C[25], Thi6_S[28], Thi6_C[28] );
FullAdder thi6fa30( Sec8_C[29], Sec9_S[27], Sec9_C[26], Thi6_S[29], Thi6_C[29] );
FullAdder thi6fa31( Sec8_C[30], Sec9_S[28], Sec9_C[27], Thi6_S[30], Thi6_C[30] );
FullAdder thi6fa32( Sec8_C[31], Sec9_S[29], Sec9_C[28], Thi6_S[31], Thi6_C[31] );
HalfAdder thi6fa33( Sec9_S[30], Sec9_C[29], Thi6_S[32], Thi6_C[32]);
HalfAdder thi6fa34( Sec9_S[31], Sec9_C[30], Thi6_S[33], Thi6_C[33]);


FullAdder thi7fa1( Sec10_C[0], Sec10_S[1], pp30[0], Thi7_S[0], Thi7_C[0] );
FullAdder thi7fa2( Sec10_C[1], Sec10_S[2], Fir11_S_[0], Thi7_S[1], Thi7_C[1] );
FullAdder thi7fa3( Sec10_C[2], Sec10_S[3], Sec11_S[0], Thi7_S[2], Thi7_C[2] );
FullAdder thi7fa4( Sec10_C[3], Sec10_S[4], Sec11_S[1], Thi7_S[3], Thi7_C[3] );
FullAdder thi7fa5( Sec10_C[4], Sec10_S[5], Sec11_S[2], Thi7_S[4], Thi7_C[4] );
FullAdder thi7fa6( Sec10_C[5], Sec10_S[6], Sec11_S[3], Thi7_S[5], Thi7_C[5] );
FullAdder thi7fa7( Sec10_C[6], Sec10_S[7], Sec11_S[4], Thi7_S[6], Thi7_C[6] );
FullAdder thi7fa8( Sec10_C[7], Sec10_S[8], Sec11_S[5], Thi7_S[7], Thi7_C[7] );
FullAdder thi7fa9( Sec10_C[8], Sec10_S[9], Sec11_S[6], Thi7_S[8], Thi7_C[8] );
FullAdder thi7fa10( Sec10_C[9], Sec10_S[10], Sec11_S[7], Thi7_S[9], Thi7_C[9] );
FullAdder thi7fa11( Sec10_C[10], Sec10_S[11], Sec11_S[8], Thi7_S[10], Thi7_C[10] );
FullAdder thi7fa12( Sec10_C[11], Sec10_S[12], Sec11_S[9], Thi7_S[11], Thi7_C[11] );
FullAdder thi7fa13( Sec10_C[12], Sec10_S[13], Sec11_S[10], Thi7_S[12], Thi7_C[12] );
FullAdder thi7fa14( Sec10_C[13], Sec10_S[14], Sec11_S[11], Thi7_S[13], Thi7_C[13] );
FullAdder thi7fa15( Sec10_C[14], Sec10_S[15], Sec11_S[12], Thi7_S[14], Thi7_C[14] );
FullAdder thi7fa16( Sec10_C[15], Sec10_S[16], Sec11_S[13], Thi7_S[15], Thi7_C[15] );
FullAdder thi7fa17( Sec10_C[16], Sec10_S[17], Sec11_S[14], Thi7_S[16], Thi7_C[16] );
FullAdder thi7fa18( Sec10_C[17], Sec10_S[18], Sec11_S[15], Thi7_S[17], Thi7_C[17] );
FullAdder thi7fa19( Sec10_C[18], Sec10_S[19], Sec11_S[16], Thi7_S[18], Thi7_C[18] );
FullAdder thi7fa20( Sec10_C[19], Sec10_S[20], Sec11_S[17], Thi7_S[19], Thi7_C[19] );
FullAdder thi7fa21( Sec10_C[20], Sec10_S[21], Sec11_S[18], Thi7_S[20], Thi7_C[20] );
FullAdder thi7fa22( Sec10_C[21], Sec10_S[22], Sec11_S[19], Thi7_S[21], Thi7_C[21] );
FullAdder thi7fa23( Sec10_C[22], Sec10_S[23], Sec11_S[20], Thi7_S[22], Thi7_C[22] );
FullAdder thi7fa24( Sec10_C[23], Sec10_S[24], Sec11_S[21], Thi7_S[23], Thi7_C[23] );
FullAdder thi7fa25( Sec10_C[24], Sec10_S[25], Sec11_S[22], Thi7_S[24], Thi7_C[24] );
FullAdder thi7fa26( Sec10_C[25], Sec10_S[26], Sec11_S[23], Thi7_S[25], Thi7_C[25] );
FullAdder thi7fa27( Sec10_C[26], Sec10_S[27], Sec11_S[24], Thi7_S[26], Thi7_C[26] );
FullAdder thi7fa28( Sec10_C[27], Sec10_S[28], Sec11_S[25], Thi7_S[27], Thi7_C[27] );
FullAdder thi7fa29( Sec10_C[28], Sec10_S[29], Sec11_S[26], Thi7_S[28], Thi7_C[28] );
FullAdder thi7fa30( Sec10_C[29], Sec10_S[30], Sec11_S[27], Thi7_S[29], Thi7_C[29] );
FullAdder thi7fa31( Sec10_C[30], Sec10_S[31], Sec11_S[28], Thi7_S[30], Thi7_C[30] );
HalfAdder thi7fa32( Sec10_C[31], Sec11_S[29], Thi7_S[31], Thi7_C[31] );



reg	[31: 0]	Thi1_S_, Thi1_C_;
reg	[33: 0]	Thi2_S_, Thi2_C_;
reg	[31: 0]	Thi3_S_, Thi3_C_;
reg	[33: 0]	Thi4_S_, Thi4_C_;
reg	[31: 0]	Thi5_S_, Thi5_C_;
reg	[33: 0]	Thi6_S_, Thi6_C_;
reg	[31: 0]	Thi7_S_, Thi7_C_;


reg done2;
reg state_done2;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Thi1_S_ <= 32'b0; Thi1_C_ <= 32'b0;
        Thi2_S_ <= 34'b0; Thi2_C_ <= 34'b0;
        Thi3_S_ <= 32'b0; Thi3_C_ <= 32'b0;
        Thi4_S_ <= 34'b0; Thi4_C_ <= 34'b0;
        Thi5_S_ <= 32'b0; Thi5_C_ <= 32'b0;
        Thi6_S_ <= 34'b0; Thi6_C_ <= 34'b0;
        Thi7_S_ <= 32'b0; Thi7_C_ <= 32'b0;
        done2 <= 1'b0;
        state_done2 <= 1'b0;
    end else begin
        case (state_done2)
            1'b0: begin
                if (done1) begin
                    Thi1_S_ <= Thi1_S; Thi1_C_ <= Thi1_C;
                    Thi2_S_ <= Thi2_S; Thi2_C_ <= Thi2_C;
                    Thi3_S_ <= Thi3_S; Thi3_C_ <= Thi3_C;
                    Thi4_S_ <= Thi4_S; Thi4_C_ <= Thi4_C;
                    Thi5_S_ <= Thi5_S; Thi5_C_ <= Thi5_C;
                    Thi6_S_ <= Thi6_S; Thi6_C_ <= Thi6_C;
                    Thi7_S_ <= Thi7_S; Thi7_C_ <= Thi7_C;
                    done2 <= 1'b1;
                    state_done2 <= 1'b1;
                end else begin
                    done2 <= 1'b0;
                end
            end
            1'b1: begin
                done2 <= 1'b0;
                if (!done1)
                    state_done2 <= 1'b0;  // Á≠âÂæÖ done1 Âèò‰∏∫ 0ÔºåÂÜçÂÖÅËÆ∏‰∏ã‰∏ÄÊ¨°ÈááÊ†?
            end
        endcase
    end
end



//===================Fourth stage===============================

wire	[31: 0]	Fou1_S_, Fou1_C_;
wire	[33: 0]	Fou2_S_, Fou2_C_;
wire	[31: 0]	Fou3_S_, Fou3_C_;
wire	[33: 0]	Fou4_S_, Fou4_C_;
wire	[31: 0]	Fou5_S_, Fou5_C_;
wire	[33: 0]	Fou6_S_, Fou6_C_;
wire	[31: 0]	Fou7_S_, Fou7_C_;


HalfAdder fou1fa1( Thi1_C_[0], Thi1_S_[1], Fou1_S_[0], Fou1_C_[0] );
HalfAdder fou1fa2( Thi1_C_[1], Thi1_S_[2], Fou1_S_[1], Fou1_C_[1] );
HalfAdder fou1fa3( Thi1_C_[2], Thi1_S_[3], Fou1_S_[2], Fou1_C_[2] );
HalfAdder fou1fa4( Thi1_C_[3], Thi1_S_[4], Fou1_S_[3], Fou1_C_[3] );
HalfAdder fou1fa5( Thi1_C_[4], Thi1_S_[5], Fou1_S_[4], Fou1_C_[4] );
HalfAdder fou1fa6( Thi1_C_[5], Thi1_S_[6], Fou1_S_[5], Fou1_C_[5] );
HalfAdder fou1fa7( Thi1_C_[6], Thi1_S_[7], Fou1_S_[6], Fou1_C_[6] );
HalfAdder fou1fa8( Thi1_C_[7], Thi1_S_[8], Fou1_S_[7], Fou1_C_[7] );
HalfAdder fou1fa9( Thi1_C_[8], Thi1_S_[9], Fou1_S_[8], Fou1_C_[8] );
HalfAdder fou1fa10( Thi1_C_[9], Thi1_S_[10], Fou1_S_[9], Fou1_C_[9] );
HalfAdder fou1fa11( Thi1_C_[10], Thi1_S_[11], Fou1_S_[10], Fou1_C_[10] );
HalfAdder fou1fa12( Thi1_C_[11], Thi1_S_[12], Fou1_S_[11], Fou1_C_[11] );
HalfAdder fou1fa13( Thi1_C_[12], Thi1_S_[13], Fou1_S_[12], Fou1_C_[12] );
HalfAdder fou1fa14( Thi1_C_[13], Thi1_S_[14], Fou1_S_[13], Fou1_C_[13] );
HalfAdder fou1fa15( Thi1_C_[14], Thi1_S_[15], Fou1_S_[14], Fou1_C_[14] );
HalfAdder fou1fa16( Thi1_C_[15], Thi1_S_[16], Fou1_S_[15], Fou1_C_[15] );
HalfAdder fou1fa17( Thi1_C_[16], Thi1_S_[17], Fou1_S_[16], Fou1_C_[16] );
HalfAdder fou1fa18( Thi1_C_[17], Thi1_S_[18], Fou1_S_[17], Fou1_C_[17] );
HalfAdder fou1fa19( Thi1_C_[18], Thi1_S_[19], Fou1_S_[18], Fou1_C_[18] );
HalfAdder fou1fa20( Thi1_C_[19], Thi1_S_[20], Fou1_S_[19], Fou1_C_[19] );
HalfAdder fou1fa21( Thi1_C_[20], Thi1_S_[21], Fou1_S_[20], Fou1_C_[20] );
HalfAdder fou1fa22( Thi1_C_[21], Thi1_S_[22], Fou1_S_[21], Fou1_C_[21] );
HalfAdder fou1fa23( Thi1_C_[22], Thi1_S_[23], Fou1_S_[22], Fou1_C_[22] );
HalfAdder fou1fa24( Thi1_C_[23], Thi1_S_[24], Fou1_S_[23], Fou1_C_[23] );
HalfAdder fou1fa25( Thi1_C_[24], Thi1_S_[25], Fou1_S_[24], Fou1_C_[24] );
HalfAdder fou1fa26( Thi1_C_[25], Thi1_S_[26], Fou1_S_[25], Fou1_C_[25] );
HalfAdder fou1fa27( Thi1_C_[26], Thi1_S_[27], Fou1_S_[26], Fou1_C_[26] );
HalfAdder fou1fa28( Thi1_C_[27], Thi1_S_[28], Fou1_S_[27], Fou1_C_[27] );
HalfAdder fou1fa29( Thi1_C_[28], Thi1_S_[29], Fou1_S_[28], Fou1_C_[28] );
HalfAdder fou1fa30( Thi1_C_[29], Thi1_S_[30], Fou1_S_[29], Fou1_C_[29] );
HalfAdder fou1fa31( Thi1_C_[30], Thi1_S_[31], Fou1_S_[30], Fou1_C_[30] );
HalfAdder fou1fa32( Thi1_C_[31], Sec2_S[30], Fou1_S_[31], Fou1_C_[31] );



HalfAdder fou2fa1( Thi2_C_[0], Thi2_S_[1], Fou2_S_[0], Fou2_C_[0] );
HalfAdder fou2fa2( Thi2_C_[1], Thi2_S_[2], Fou2_S_[1], Fou2_C_[1] );
HalfAdder fou2fa3( Thi2_C_[2], Thi2_S_[3], Fou2_S_[2], Fou2_C_[2] );
HalfAdder fou2fa4( Thi2_C_[3], Thi2_S_[4], Fou2_S_[3], Fou2_C_[3] );
HalfAdder fou2fa5( Thi2_C_[4], Thi2_S_[5], Fou2_S_[4], Fou2_C_[4] );
HalfAdder fou2fa6( Thi2_C_[5], Thi2_S_[6], Fou2_S_[5], Fou2_C_[5] );
HalfAdder fou2fa7( Thi2_C_[6], Thi2_S_[7], Fou2_S_[6], Fou2_C_[6] );
HalfAdder fou2fa8( Thi2_C_[7], Thi2_S_[8], Fou2_S_[7], Fou2_C_[7] );
HalfAdder fou2fa9( Thi2_C_[8], Thi2_S_[9], Fou2_S_[8], Fou2_C_[8] );
HalfAdder fou2fa10( Thi2_C_[9], Thi2_S_[10], Fou2_S_[9], Fou2_C_[9] );
HalfAdder fou2fa11( Thi2_C_[10], Thi2_S_[11], Fou2_S_[10], Fou2_C_[10] );
HalfAdder fou2fa12( Thi2_C_[11], Thi2_S_[12], Fou2_S_[11], Fou2_C_[11] );
HalfAdder fou2fa13( Thi2_C_[12], Thi2_S_[13], Fou2_S_[12], Fou2_C_[12] );
HalfAdder fou2fa14( Thi2_C_[13], Thi2_S_[14], Fou2_S_[13], Fou2_C_[13] );
HalfAdder fou2fa15( Thi2_C_[14], Thi2_S_[15], Fou2_S_[14], Fou2_C_[14] );
HalfAdder fou2fa16( Thi2_C_[15], Thi2_S_[16], Fou2_S_[15], Fou2_C_[15] );
HalfAdder fou2fa17( Thi2_C_[16], Thi2_S_[17], Fou2_S_[16], Fou2_C_[16] );
HalfAdder fou2fa18( Thi2_C_[17], Thi2_S_[18], Fou2_S_[17], Fou2_C_[17] );
HalfAdder fou2fa19( Thi2_C_[18], Thi2_S_[19], Fou2_S_[18], Fou2_C_[18] );
HalfAdder fou2fa20( Thi2_C_[19], Thi2_S_[20], Fou2_S_[19], Fou2_C_[19] );
HalfAdder fou2fa21( Thi2_C_[20], Thi2_S_[21], Fou2_S_[20], Fou2_C_[20] );
HalfAdder fou2fa22( Thi2_C_[21], Thi2_S_[22], Fou2_S_[21], Fou2_C_[21] );
HalfAdder fou2fa23( Thi2_C_[22], Thi2_S_[23], Fou2_S_[22], Fou2_C_[22] );
HalfAdder fou2fa24( Thi2_C_[23], Thi2_S_[24], Fou2_S_[23], Fou2_C_[23] );
HalfAdder fou2fa25( Thi2_C_[24], Thi2_S_[25], Fou2_S_[24], Fou2_C_[24] );
HalfAdder fou2fa26( Thi2_C_[25], Thi2_S_[26], Fou2_S_[25], Fou2_C_[25] );
HalfAdder fou2fa27( Thi2_C_[26], Thi2_S_[27], Fou2_S_[26], Fou2_C_[26] );
HalfAdder fou2fa28( Thi2_C_[27], Thi2_S_[28], Fou2_S_[27], Fou2_C_[27] );
HalfAdder fou2fa29( Thi2_C_[28], Thi2_S_[29], Fou2_S_[28], Fou2_C_[28] );
HalfAdder fou2fa30( Thi2_C_[29], Thi2_S_[30], Fou2_S_[29], Fou2_C_[29] );
HalfAdder fou2fa31( Thi2_C_[30], Thi2_S_[31], Fou2_S_[30], Fou2_C_[30] );
HalfAdder fou2fa32( Thi2_C_[31], Thi2_S_[32], Fou2_S_[31], Fou2_C_[31] );
HalfAdder fou2fa33( Thi2_C_[32], Thi2_S_[33], Fou2_S_[32], Fou2_C_[32] );
HalfAdder fou2fa34( Thi2_C_[33], Sec3_C[31], Fou2_S_[33], Fou2_C_[33] );



HalfAdder fou3fa1( Thi3_C_[0], Thi3_S_[1], Fou3_S_[0], Fou3_C_[0] );
HalfAdder fou3fa2( Thi3_C_[1], Thi3_S_[2], Fou3_S_[1], Fou3_C_[1] );
HalfAdder fou3fa3( Thi3_C_[2], Thi3_S_[3], Fou3_S_[2], Fou3_C_[2] );
HalfAdder fou3fa4( Thi3_C_[3], Thi3_S_[4], Fou3_S_[3], Fou3_C_[3] );
HalfAdder fou3fa5( Thi3_C_[4], Thi3_S_[5], Fou3_S_[4], Fou3_C_[4] );
HalfAdder fou3fa6( Thi3_C_[5], Thi3_S_[6], Fou3_S_[5], Fou3_C_[5] );
HalfAdder fou3fa7( Thi3_C_[6], Thi3_S_[7], Fou3_S_[6], Fou3_C_[6] );
HalfAdder fou3fa8( Thi3_C_[7], Thi3_S_[8], Fou3_S_[7], Fou3_C_[7] );
HalfAdder fou3fa9( Thi3_C_[8], Thi3_S_[9], Fou3_S_[8], Fou3_C_[8] );
HalfAdder fou3fa10( Thi3_C_[9], Thi3_S_[10], Fou3_S_[9], Fou3_C_[9] );
HalfAdder fou3fa11( Thi3_C_[10], Thi3_S_[11], Fou3_S_[10], Fou3_C_[10] );
HalfAdder fou3fa12( Thi3_C_[11], Thi3_S_[12], Fou3_S_[11], Fou3_C_[11] );
HalfAdder fou3fa13( Thi3_C_[12], Thi3_S_[13], Fou3_S_[12], Fou3_C_[12] );
HalfAdder fou3fa14( Thi3_C_[13], Thi3_S_[14], Fou3_S_[13], Fou3_C_[13] );
HalfAdder fou3fa15( Thi3_C_[14], Thi3_S_[15], Fou3_S_[14], Fou3_C_[14] );
HalfAdder fou3fa16( Thi3_C_[15], Thi3_S_[16], Fou3_S_[15], Fou3_C_[15] );
HalfAdder fou3fa17( Thi3_C_[16], Thi3_S_[17], Fou3_S_[16], Fou3_C_[16] );
HalfAdder fou3fa18( Thi3_C_[17], Thi3_S_[18], Fou3_S_[17], Fou3_C_[17] );
HalfAdder fou3fa19( Thi3_C_[18], Thi3_S_[19], Fou3_S_[18], Fou3_C_[18] );
HalfAdder fou3fa20( Thi3_C_[19], Thi3_S_[20], Fou3_S_[19], Fou3_C_[19] );
HalfAdder fou3fa21( Thi3_C_[20], Thi3_S_[21], Fou3_S_[20], Fou3_C_[20] );
HalfAdder fou3fa22( Thi3_C_[21], Thi3_S_[22], Fou3_S_[21], Fou3_C_[21] );
HalfAdder fou3fa23( Thi3_C_[22], Thi3_S_[23], Fou3_S_[22], Fou3_C_[22] );
HalfAdder fou3fa24( Thi3_C_[23], Thi3_S_[24], Fou3_S_[23], Fou3_C_[23] );
HalfAdder fou3fa25( Thi3_C_[24], Thi3_S_[25], Fou3_S_[24], Fou3_C_[24] );
HalfAdder fou3fa26( Thi3_C_[25], Thi3_S_[26], Fou3_S_[25], Fou3_C_[25] );
HalfAdder fou3fa27( Thi3_C_[26], Thi3_S_[27], Fou3_S_[26], Fou3_C_[26] );
HalfAdder fou3fa28( Thi3_C_[27], Thi3_S_[28], Fou3_S_[27], Fou3_C_[27] );
HalfAdder fou3fa29( Thi3_C_[28], Thi3_S_[29], Fou3_S_[28], Fou3_C_[28] );
HalfAdder fou3fa30( Thi3_C_[29], Thi3_S_[30], Fou3_S_[29], Fou3_C_[29] );
HalfAdder fou3fa31( Thi3_C_[30], Thi3_S_[31], Fou3_S_[30], Fou3_C_[30] );
HalfAdder fou3fa32( Thi3_C_[31], Sec5_S[30], Fou3_S_[31], Fou3_C_[31] );


HalfAdder fou4fa1( Thi4_C_[0], Thi4_S_[1], Fou4_S_[0], Fou4_C_[0] );
HalfAdder fou4fa2( Thi4_C_[1], Thi4_S_[2], Fou4_S_[1], Fou4_C_[1] );
HalfAdder fou4fa3( Thi4_C_[2], Thi4_S_[3], Fou4_S_[2], Fou4_C_[2] );
HalfAdder fou4fa4( Thi4_C_[3], Thi4_S_[4], Fou4_S_[3], Fou4_C_[3] );
HalfAdder fou4fa5( Thi4_C_[4], Thi4_S_[5], Fou4_S_[4], Fou4_C_[4] );
HalfAdder fou4fa6( Thi4_C_[5], Thi4_S_[6], Fou4_S_[5], Fou4_C_[5] );
HalfAdder fou4fa7( Thi4_C_[6], Thi4_S_[7], Fou4_S_[6], Fou4_C_[6] );
HalfAdder fou4fa8( Thi4_C_[7], Thi4_S_[8], Fou4_S_[7], Fou4_C_[7] );
HalfAdder fou4fa9( Thi4_C_[8], Thi4_S_[9], Fou4_S_[8], Fou4_C_[8] );
HalfAdder fou4fa10( Thi4_C_[9], Thi4_S_[10], Fou4_S_[9], Fou4_C_[9] );
HalfAdder fou4fa11( Thi4_C_[10], Thi4_S_[11], Fou4_S_[10], Fou4_C_[10] );
HalfAdder fou4fa12( Thi4_C_[11], Thi4_S_[12], Fou4_S_[11], Fou4_C_[11] );
HalfAdder fou4fa13( Thi4_C_[12], Thi4_S_[13], Fou4_S_[12], Fou4_C_[12] );
HalfAdder fou4fa14( Thi4_C_[13], Thi4_S_[14], Fou4_S_[13], Fou4_C_[13] );
HalfAdder fou4fa15( Thi4_C_[14], Thi4_S_[15], Fou4_S_[14], Fou4_C_[14] );
HalfAdder fou4fa16( Thi4_C_[15], Thi4_S_[16], Fou4_S_[15], Fou4_C_[15] );
HalfAdder fou4fa17( Thi4_C_[16], Thi4_S_[17], Fou4_S_[16], Fou4_C_[16] );
HalfAdder fou4fa18( Thi4_C_[17], Thi4_S_[18], Fou4_S_[17], Fou4_C_[17] );
HalfAdder fou4fa19( Thi4_C_[18], Thi4_S_[19], Fou4_S_[18], Fou4_C_[18] );
HalfAdder fou4fa20( Thi4_C_[19], Thi4_S_[20], Fou4_S_[19], Fou4_C_[19] );
HalfAdder fou4fa21( Thi4_C_[20], Thi4_S_[21], Fou4_S_[20], Fou4_C_[20] );
HalfAdder fou4fa22( Thi4_C_[21], Thi4_S_[22], Fou4_S_[21], Fou4_C_[21] );
HalfAdder fou4fa23( Thi4_C_[22], Thi4_S_[23], Fou4_S_[22], Fou4_C_[22] );
HalfAdder fou4fa24( Thi4_C_[23], Thi4_S_[24], Fou4_S_[23], Fou4_C_[23] );
HalfAdder fou4fa25( Thi4_C_[24], Thi4_S_[25], Fou4_S_[24], Fou4_C_[24] );
HalfAdder fou4fa26( Thi4_C_[25], Thi4_S_[26], Fou4_S_[25], Fou4_C_[25] );
HalfAdder fou4fa27( Thi4_C_[26], Thi4_S_[27], Fou4_S_[26], Fou4_C_[26] );
HalfAdder fou4fa28( Thi4_C_[27], Thi4_S_[28], Fou4_S_[27], Fou4_C_[27] );
HalfAdder fou4fa29( Thi4_C_[28], Thi4_S_[29], Fou4_S_[28], Fou4_C_[28] );
HalfAdder fou4fa30( Thi4_C_[29], Thi4_S_[30], Fou4_S_[29], Fou4_C_[29] );
HalfAdder fou4fa31( Thi4_C_[30], Thi4_S_[31], Fou4_S_[30], Fou4_C_[30] );
HalfAdder fou4fa32( Thi4_C_[31], Thi4_S_[32], Fou4_S_[31], Fou4_C_[31] );
HalfAdder fou4fa33( Thi4_C_[32], Thi4_S_[33], Fou4_S_[32], Fou4_C_[32] );
HalfAdder fou4fa34( Thi4_C_[33], Sec6_C[31], Fou4_S_[33], Fou4_C_[33] );

HalfAdder fou5fa1( Thi5_C_[0], Thi5_S_[1], Fou5_S_[0], Fou5_C_[0] );
HalfAdder fou5fa2( Thi5_C_[1], Thi5_S_[2], Fou5_S_[1], Fou5_C_[1] );
HalfAdder fou5fa3( Thi5_C_[2], Thi5_S_[3], Fou5_S_[2], Fou5_C_[2] );
HalfAdder fou5fa4( Thi5_C_[3], Thi5_S_[4], Fou5_S_[3], Fou5_C_[3] );
HalfAdder fou5fa5( Thi5_C_[4], Thi5_S_[5], Fou5_S_[4], Fou5_C_[4] );
HalfAdder fou5fa6( Thi5_C_[5], Thi5_S_[6], Fou5_S_[5], Fou5_C_[5] );
HalfAdder fou5fa7( Thi5_C_[6], Thi5_S_[7], Fou5_S_[6], Fou5_C_[6] );
HalfAdder fou5fa8( Thi5_C_[7], Thi5_S_[8], Fou5_S_[7], Fou5_C_[7] );
HalfAdder fou5fa9( Thi5_C_[8], Thi5_S_[9], Fou5_S_[8], Fou5_C_[8] );
HalfAdder fou5fa10( Thi5_C_[9], Thi5_S_[10], Fou5_S_[9], Fou5_C_[9] );
HalfAdder fou5fa11( Thi5_C_[10], Thi5_S_[11], Fou5_S_[10], Fou5_C_[10] );
HalfAdder fou5fa12( Thi5_C_[11], Thi5_S_[12], Fou5_S_[11], Fou5_C_[11] );
HalfAdder fou5fa13( Thi5_C_[12], Thi5_S_[13], Fou5_S_[12], Fou5_C_[12] );
HalfAdder fou5fa14( Thi5_C_[13], Thi5_S_[14], Fou5_S_[13], Fou5_C_[13] );
HalfAdder fou5fa15( Thi5_C_[14], Thi5_S_[15], Fou5_S_[14], Fou5_C_[14] );
HalfAdder fou5fa16( Thi5_C_[15], Thi5_S_[16], Fou5_S_[15], Fou5_C_[15] );
HalfAdder fou5fa17( Thi5_C_[16], Thi5_S_[17], Fou5_S_[16], Fou5_C_[16] );
HalfAdder fou5fa18( Thi5_C_[17], Thi5_S_[18], Fou5_S_[17], Fou5_C_[17] );
HalfAdder fou5fa19( Thi5_C_[18], Thi5_S_[19], Fou5_S_[18], Fou5_C_[18] );
HalfAdder fou5fa20( Thi5_C_[19], Thi5_S_[20], Fou5_S_[19], Fou5_C_[19] );
HalfAdder fou5fa21( Thi5_C_[20], Thi5_S_[21], Fou5_S_[20], Fou5_C_[20] );
HalfAdder fou5fa22( Thi5_C_[21], Thi5_S_[22], Fou5_S_[21], Fou5_C_[21] );
HalfAdder fou5fa23( Thi5_C_[22], Thi5_S_[23], Fou5_S_[22], Fou5_C_[22] );
HalfAdder fou5fa24( Thi5_C_[23], Thi5_S_[24], Fou5_S_[23], Fou5_C_[23] );
HalfAdder fou5fa25( Thi5_C_[24], Thi5_S_[25], Fou5_S_[24], Fou5_C_[24] );
HalfAdder fou5fa26( Thi5_C_[25], Thi5_S_[26], Fou5_S_[25], Fou5_C_[25] );
HalfAdder fou5fa27( Thi5_C_[26], Thi5_S_[27], Fou5_S_[26], Fou5_C_[26] );
HalfAdder fou5fa28( Thi5_C_[27], Thi5_S_[28], Fou5_S_[27], Fou5_C_[27] );
HalfAdder fou5fa29( Thi5_C_[28], Thi5_S_[29], Fou5_S_[28], Fou5_C_[28] );
HalfAdder fou5fa30( Thi5_C_[29], Thi5_S_[30], Fou5_S_[29], Fou5_C_[29] );
HalfAdder fou5fa31( Thi5_C_[30], Thi5_S_[31], Fou5_S_[30], Fou5_C_[30] );
HalfAdder fou5fa32( Thi5_C_[31], Sec8_S[30], Fou5_S_[31], Fou5_C_[31] );


HalfAdder fou6fa1( Thi6_C_[0], Thi6_S_[1], Fou6_S_[0], Fou6_C_[0] );
HalfAdder fou6fa2( Thi6_C_[1], Thi6_S_[2], Fou6_S_[1], Fou6_C_[1] );
HalfAdder fou6fa3( Thi6_C_[2], Thi6_S_[3], Fou6_S_[2], Fou6_C_[2] );
HalfAdder fou6fa4( Thi6_C_[3], Thi6_S_[4], Fou6_S_[3], Fou6_C_[3] );
HalfAdder fou6fa5( Thi6_C_[4], Thi6_S_[5], Fou6_S_[4], Fou6_C_[4] );
HalfAdder fou6fa6( Thi6_C_[5], Thi6_S_[6], Fou6_S_[5], Fou6_C_[5] );
HalfAdder fou6fa7( Thi6_C_[6], Thi6_S_[7], Fou6_S_[6], Fou6_C_[6] );
HalfAdder fou6fa8( Thi6_C_[7], Thi6_S_[8], Fou6_S_[7], Fou6_C_[7] );
HalfAdder fou6fa9( Thi6_C_[8], Thi6_S_[9], Fou6_S_[8], Fou6_C_[8] );
HalfAdder fou6fa10( Thi6_C_[9], Thi6_S_[10], Fou6_S_[9], Fou6_C_[9] );
HalfAdder fou6fa11( Thi6_C_[10], Thi6_S_[11], Fou6_S_[10], Fou6_C_[10] );
HalfAdder fou6fa12( Thi6_C_[11], Thi6_S_[12], Fou6_S_[11], Fou6_C_[11] );
HalfAdder fou6fa13( Thi6_C_[12], Thi6_S_[13], Fou6_S_[12], Fou6_C_[12] );
HalfAdder fou6fa14( Thi6_C_[13], Thi6_S_[14], Fou6_S_[13], Fou6_C_[13] );
HalfAdder fou6fa15( Thi6_C_[14], Thi6_S_[15], Fou6_S_[14], Fou6_C_[14] );
HalfAdder fou6fa16( Thi6_C_[15], Thi6_S_[16], Fou6_S_[15], Fou6_C_[15] );
HalfAdder fou6fa17( Thi6_C_[16], Thi6_S_[17], Fou6_S_[16], Fou6_C_[16] );
HalfAdder fou6fa18( Thi6_C_[17], Thi6_S_[18], Fou6_S_[17], Fou6_C_[17] );
HalfAdder fou6fa19( Thi6_C_[18], Thi6_S_[19], Fou6_S_[18], Fou6_C_[18] );
HalfAdder fou6fa20( Thi6_C_[19], Thi6_S_[20], Fou6_S_[19], Fou6_C_[19] );
HalfAdder fou6fa21( Thi6_C_[20], Thi6_S_[21], Fou6_S_[20], Fou6_C_[20] );
HalfAdder fou6fa22( Thi6_C_[21], Thi6_S_[22], Fou6_S_[21], Fou6_C_[21] );
HalfAdder fou6fa23( Thi6_C_[22], Thi6_S_[23], Fou6_S_[22], Fou6_C_[22] );
HalfAdder fou6fa24( Thi6_C_[23], Thi6_S_[24], Fou6_S_[23], Fou6_C_[23] );
HalfAdder fou6fa25( Thi6_C_[24], Thi6_S_[25], Fou6_S_[24], Fou6_C_[24] );
HalfAdder fou6fa26( Thi6_C_[25], Thi6_S_[26], Fou6_S_[25], Fou6_C_[25] );
HalfAdder fou6fa27( Thi6_C_[26], Thi6_S_[27], Fou6_S_[26], Fou6_C_[26] );
HalfAdder fou6fa28( Thi6_C_[27], Thi6_S_[28], Fou6_S_[27], Fou6_C_[27] );
HalfAdder fou6fa29( Thi6_C_[28], Thi6_S_[29], Fou6_S_[28], Fou6_C_[28] );
HalfAdder fou6fa30( Thi6_C_[29], Thi6_S_[30], Fou6_S_[29], Fou6_C_[29] );
HalfAdder fou6fa31( Thi6_C_[30], Thi6_S_[31], Fou6_S_[30], Fou6_C_[30] );
HalfAdder fou6fa32( Thi6_C_[31], Thi6_S_[32], Fou6_S_[31], Fou6_C_[31] );
HalfAdder fou6fa33( Thi6_C_[32], Thi6_S_[33], Fou6_S_[32], Fou6_C_[32] );
HalfAdder fou6fa34( Thi6_C_[33], Sec9_C[31], Fou6_S_[33], Fou6_C_[33] );

HalfAdder fou7fa1( Thi7_C_[0], Thi7_S_[1], Fou7_S_[0], Fou7_C_[0] );
HalfAdder fou7fa2( Thi7_C_[1], Thi7_S_[2], Fou7_S_[1], Fou7_C_[1] );
HalfAdder fou7fa3( Thi7_C_[2], Thi7_S_[3], Fou7_S_[2], Fou7_C_[2] );
HalfAdder fou7fa4( Thi7_C_[3], Thi7_S_[4], Fou7_S_[3], Fou7_C_[3] );
HalfAdder fou7fa5( Thi7_C_[4], Thi7_S_[5], Fou7_S_[4], Fou7_C_[4] );
HalfAdder fou7fa6( Thi7_C_[5], Thi7_S_[6], Fou7_S_[5], Fou7_C_[5] );
HalfAdder fou7fa7( Thi7_C_[6], Thi7_S_[7], Fou7_S_[6], Fou7_C_[6] );
HalfAdder fou7fa8( Thi7_C_[7], Thi7_S_[8], Fou7_S_[7], Fou7_C_[7] );
HalfAdder fou7fa9( Thi7_C_[8], Thi7_S_[9], Fou7_S_[8], Fou7_C_[8] );
HalfAdder fou7fa10( Thi7_C_[9], Thi7_S_[10], Fou7_S_[9], Fou7_C_[9] );
HalfAdder fou7fa11( Thi7_C_[10], Thi7_S_[11], Fou7_S_[10], Fou7_C_[10] );
HalfAdder fou7fa12( Thi7_C_[11], Thi7_S_[12], Fou7_S_[11], Fou7_C_[11] );
HalfAdder fou7fa13( Thi7_C_[12], Thi7_S_[13], Fou7_S_[12], Fou7_C_[12] );
HalfAdder fou7fa14( Thi7_C_[13], Thi7_S_[14], Fou7_S_[13], Fou7_C_[13] );
HalfAdder fou7fa15( Thi7_C_[14], Thi7_S_[15], Fou7_S_[14], Fou7_C_[14] );
HalfAdder fou7fa16( Thi7_C_[15], Thi7_S_[16], Fou7_S_[15], Fou7_C_[15] );
HalfAdder fou7fa17( Thi7_C_[16], Thi7_S_[17], Fou7_S_[16], Fou7_C_[16] );
HalfAdder fou7fa18( Thi7_C_[17], Thi7_S_[18], Fou7_S_[17], Fou7_C_[17] );
HalfAdder fou7fa19( Thi7_C_[18], Thi7_S_[19], Fou7_S_[18], Fou7_C_[18] );
HalfAdder fou7fa20( Thi7_C_[19], Thi7_S_[20], Fou7_S_[19], Fou7_C_[19] );
HalfAdder fou7fa21( Thi7_C_[20], Thi7_S_[21], Fou7_S_[20], Fou7_C_[20] );
HalfAdder fou7fa22( Thi7_C_[21], Thi7_S_[22], Fou7_S_[21], Fou7_C_[21] );
HalfAdder fou7fa23( Thi7_C_[22], Thi7_S_[23], Fou7_S_[22], Fou7_C_[22] );
HalfAdder fou7fa24( Thi7_C_[23], Thi7_S_[24], Fou7_S_[23], Fou7_C_[23] );
HalfAdder fou7fa25( Thi7_C_[24], Thi7_S_[25], Fou7_S_[24], Fou7_C_[24] );
HalfAdder fou7fa26( Thi7_C_[25], Thi7_S_[26], Fou7_S_[25], Fou7_C_[25] );
HalfAdder fou7fa27( Thi7_C_[26], Thi7_S_[27], Fou7_S_[26], Fou7_C_[26] );
HalfAdder fou7fa28( Thi7_C_[27], Thi7_S_[28], Fou7_S_[27], Fou7_C_[27] );
HalfAdder fou7fa29( Thi7_C_[28], Thi7_S_[29], Fou7_S_[28], Fou7_C_[28] );
HalfAdder fou7fa30( Thi7_C_[29], Thi7_S_[30], Fou7_S_[29], Fou7_C_[29] );
HalfAdder fou7fa31( Thi7_C_[30], Thi7_S_[31], Fou7_S_[30], Fou7_C_[30] );
HalfAdder fou7fa32( Thi7_C_[31], Sec11_S[30], Fou7_S_[31], Fou7_C_[31] );


reg	[31: 0]	Fou1_S, Fou1_C;
reg	[33: 0]	Fou2_S, Fou2_C;
reg	[31: 0]	Fou3_S, Fou3_C;
reg	[33: 0]	Fou4_S, Fou4_C;
reg	[31: 0]	Fou5_S, Fou5_C;
reg	[33: 0]	Fou6_S, Fou6_C;
reg	[31: 0]	Fou7_S, Fou7_C;

reg done3;
reg state_done3;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Fou1_S <= 32'b0; Fou1_C <= 32'b0;
        Fou2_S <= 34'b0; Fou2_C <= 34'b0;
        Fou3_S <= 32'b0; Fou3_C <= 32'b0;
        Fou4_S <= 34'b0; Fou4_C <= 34'b0;
        Fou5_S <= 32'b0; Fou5_C <= 32'b0;
        Fou6_S <= 34'b0; Fou6_C <= 34'b0;
        Fou7_S <= 32'b0; Fou7_C <= 32'b0;
        done3 <= 1'b0;
        state_done3 <= 1'b0;
    end else begin
        case (state_done3)
            1'b0: begin
                if (done2) begin
                    Fou1_S <= Fou1_S_; Fou1_C <= Fou1_C_;
                    Fou2_S <= Fou2_S_; Fou2_C <= Fou2_C_;
                    Fou3_S <= Fou3_S_; Fou3_C <= Fou3_C_;
                    Fou4_S <= Fou4_S_; Fou4_C <= Fou4_C_;
                    Fou5_S <= Fou5_S_; Fou5_C <= Fou5_C_;
                    Fou6_S <= Fou6_S_; Fou6_C <= Fou6_C_;
                    Fou7_S <= Fou7_S_; Fou7_C <= Fou7_C_;
                    done3 <= 1'b1;
                    state_done3 <= 1'b1;
                end else begin
                    done3 <= 1'b0;
                end
            end
            1'b1: begin
                done3 <= 1'b0;
                if (!done2)
                    state_done3 <= 1'b0;
            end
        endcase
    end
end



//===================Fifth stage===============================

wire	[31: 0]	Fif1_S, Fif1_C;
wire	[36: 0]	Fif2_S, Fif2_C;
wire	[33: 0]	Fif3_S, Fif3_C;
wire	[34: 0]	Fif4_S, Fif4_C;
wire	[31: 0]	Fif5_S, Fif5_C;




HalfAdder fif1fa1( Fou1_C[0], Fou1_S[1], Fif1_S[0], Fif1_C[0] );
FullAdder fif1fa2( Fou1_C[1], Fou1_S[2], Thi2_S_[0], Fif1_S[1], Fif1_C[1] );
FullAdder fif1fa3( Fou1_C[2], Fou1_S[3], Fou2_S[0], Fif1_S[2], Fif1_C[2] );
FullAdder fif1fa4( Fou1_C[3], Fou1_S[4], Fou2_S[1], Fif1_S[3], Fif1_C[3] );
FullAdder fif1fa5( Fou1_C[4], Fou1_S[5], Fou2_S[2], Fif1_S[4], Fif1_C[4] );
FullAdder fif1fa6( Fou1_C[5], Fou1_S[6], Fou2_S[3], Fif1_S[5], Fif1_C[5] );
FullAdder fif1fa7( Fou1_C[6], Fou1_S[7], Fou2_S[4], Fif1_S[6], Fif1_C[6] );
FullAdder fif1fa8( Fou1_C[7], Fou1_S[8], Fou2_S[5], Fif1_S[7], Fif1_C[7] );
FullAdder fif1fa9( Fou1_C[8], Fou1_S[9], Fou2_S[6], Fif1_S[8], Fif1_C[8] );
FullAdder fif1fa10( Fou1_C[9], Fou1_S[10], Fou2_S[7], Fif1_S[9], Fif1_C[9] );
FullAdder fif1fa11( Fou1_C[10], Fou1_S[11], Fou2_S[8], Fif1_S[10], Fif1_C[10] );
FullAdder fif1fa12( Fou1_C[11], Fou1_S[12], Fou2_S[9], Fif1_S[11], Fif1_C[11] );
FullAdder fif1fa13( Fou1_C[12], Fou1_S[13], Fou2_S[10], Fif1_S[12], Fif1_C[12] );
FullAdder fif1fa14( Fou1_C[13], Fou1_S[14], Fou2_S[11], Fif1_S[13], Fif1_C[13] );
FullAdder fif1fa15( Fou1_C[14], Fou1_S[15], Fou2_S[12], Fif1_S[14], Fif1_C[14] );
FullAdder fif1fa16( Fou1_C[15], Fou1_S[16], Fou2_S[13], Fif1_S[15], Fif1_C[15] );
FullAdder fif1fa17( Fou1_C[16], Fou1_S[17], Fou2_S[14], Fif1_S[16], Fif1_C[16] );
FullAdder fif1fa18( Fou1_C[17], Fou1_S[18], Fou2_S[15], Fif1_S[17], Fif1_C[17] );
FullAdder fif1fa19( Fou1_C[18], Fou1_S[19], Fou2_S[16], Fif1_S[18], Fif1_C[18] );
FullAdder fif1fa20( Fou1_C[19], Fou1_S[20], Fou2_S[17], Fif1_S[19], Fif1_C[19] );
FullAdder fif1fa21( Fou1_C[20], Fou1_S[21], Fou2_S[18], Fif1_S[20], Fif1_C[20] );
FullAdder fif1fa22( Fou1_C[21], Fou1_S[22], Fou2_S[19], Fif1_S[21], Fif1_C[21] );
FullAdder fif1fa23( Fou1_C[22], Fou1_S[23], Fou2_S[20], Fif1_S[22], Fif1_C[22] );
FullAdder fif1fa24( Fou1_C[23], Fou1_S[24], Fou2_S[21], Fif1_S[23], Fif1_C[23] );
FullAdder fif1fa25( Fou1_C[24], Fou1_S[25], Fou2_S[22], Fif1_S[24], Fif1_C[24] );
FullAdder fif1fa26( Fou1_C[25], Fou1_S[26], Fou2_S[23], Fif1_S[25], Fif1_C[25] );
FullAdder fif1fa27( Fou1_C[26], Fou1_S[27], Fou2_S[24], Fif1_S[26], Fif1_C[26] );
FullAdder fif1fa28( Fou1_C[27], Fou1_S[28], Fou2_S[25], Fif1_S[27], Fif1_C[27] );
FullAdder fif1fa29( Fou1_C[28], Fou1_S[29], Fou2_S[26], Fif1_S[28], Fif1_C[28] );
FullAdder fif1fa30( Fou1_C[29], Fou1_S[30], Fou2_S[27], Fif1_S[29], Fif1_C[29] );
FullAdder fif1fa31( Fou1_C[30], Fou1_S[31], Fou2_S[28], Fif1_S[30], Fif1_C[30] );
FullAdder fif1fa32( Fou1_C[31], Sec2_S[31], Fou2_S[29], Fif1_S[31], Fif1_C[31] );

HalfAdder fif2fa1( pp9[0], Fou2_C[1], Fif2_S[0], Fif2_C[0] );
HalfAdder fif2fa2( Fir4_S_[0], Fou2_C[2], Fif2_S[1], Fif2_C[1] );
HalfAdder fif2fa3( Sec4_S[0], Fou2_C[3], Fif2_S[2], Fif2_C[2] );
HalfAdder fif2fa4(Thi3_S_[0], Fou2_C[4], Fif2_S[3], Fif2_C[3] );
HalfAdder fif2fa5( Fou3_S[0], Fou2_C[5], Fif2_S[4], Fif2_C[4] );
FullAdder fif2fa6( Fou3_S[1], Fou2_C[6], Fou3_C[0], Fif2_S[5], Fif2_C[5] );
FullAdder fif2fa7( Fou3_S[2], Fou2_C[7], Fou3_C[1], Fif2_S[6], Fif2_C[6] );
FullAdder fif2fa8( Fou3_S[3], Fou2_C[8], Fou3_C[2], Fif2_S[7], Fif2_C[7] );
FullAdder fif2fa9( Fou3_S[4], Fou2_C[9], Fou3_C[3], Fif2_S[8], Fif2_C[8] );
FullAdder fif2fa10( Fou3_S[5], Fou2_C[10], Fou3_C[4], Fif2_S[9], Fif2_C[9] );
FullAdder fif2fa11( Fou3_S[6], Fou2_C[11], Fou3_C[5], Fif2_S[10], Fif2_C[10] );
FullAdder fif2fa12( Fou3_S[7], Fou2_C[12], Fou3_C[6], Fif2_S[11], Fif2_C[11] );
FullAdder fif2fa13( Fou3_S[8], Fou2_C[13], Fou3_C[7], Fif2_S[12], Fif2_C[12] );
FullAdder fif2fa14( Fou3_S[9], Fou2_C[14], Fou3_C[8], Fif2_S[13], Fif2_C[13] );
FullAdder fif2fa15( Fou3_S[10], Fou2_C[15], Fou3_C[9], Fif2_S[14], Fif2_C[14] );
FullAdder fif2fa16( Fou3_S[11], Fou2_C[16], Fou3_C[10], Fif2_S[15], Fif2_C[15] );
FullAdder fif2fa17( Fou3_S[12], Fou2_C[17], Fou3_C[11], Fif2_S[16], Fif2_C[16] );
FullAdder fif2fa18( Fou3_S[13], Fou2_C[18], Fou3_C[12], Fif2_S[17], Fif2_C[17] );
FullAdder fif2fa19( Fou3_S[14], Fou2_C[19], Fou3_C[13], Fif2_S[18], Fif2_C[18] );
FullAdder fif2fa20( Fou3_S[15], Fou2_C[20], Fou3_C[14], Fif2_S[19], Fif2_C[19] );
FullAdder fif2fa21( Fou3_S[16], Fou2_C[21], Fou3_C[15], Fif2_S[20], Fif2_C[20] );
FullAdder fif2fa22( Fou3_S[17], Fou2_C[22], Fou3_C[16], Fif2_S[21], Fif2_C[21] );
FullAdder fif2fa23( Fou3_S[18], Fou2_C[23], Fou3_C[17], Fif2_S[22], Fif2_C[22] );
FullAdder fif2fa24( Fou3_S[19], Fou2_C[24], Fou3_C[18], Fif2_S[23], Fif2_C[23] );
FullAdder fif2fa25( Fou3_S[20], Fou2_C[25], Fou3_C[19], Fif2_S[24], Fif2_C[24] );
FullAdder fif2fa26( Fou3_S[21], Fou2_C[26], Fou3_C[20], Fif2_S[25], Fif2_C[25] );
FullAdder fif2fa27( Fou3_S[22], Fou2_C[27], Fou3_C[21], Fif2_S[26], Fif2_C[26] );
FullAdder fif2fa28( Fou3_S[23], Fou2_C[28], Fou3_C[22], Fif2_S[27], Fif2_C[27] );
FullAdder fif2fa29( Fou3_S[24], Fou2_C[29], Fou3_C[23], Fif2_S[28], Fif2_C[28] );
FullAdder fif2fa30( Fou3_S[25], Fou2_C[30], Fou3_C[24], Fif2_S[29], Fif2_C[29] );
FullAdder fif2fa31( Fou3_S[26], Fou2_C[31], Fou3_C[25], Fif2_S[30], Fif2_C[30] );
FullAdder fif2fa32( Fou3_S[27], Fou2_C[32], Fou3_C[26], Fif2_S[31], Fif2_C[31] );
FullAdder fif2fa33( Fou3_S[28], Fou2_C[33], Fou3_C[27], Fif2_S[32], Fif2_C[32] );
HalfAdder fif2fa34( Fou3_S[29], Fou3_C[28], Fif2_S[33], Fif2_C[33] );
HalfAdder fif2fa35( Fou3_S[30], Fou3_C[29], Fif2_S[34], Fif2_C[34] );
HalfAdder fif2fa36( Fou3_S[31], Fou3_C[30], Fif2_S[35], Fif2_C[35] );
HalfAdder fif2fa37( Sec5_S[31], Fou3_C[31], Fif2_S[36], Fif2_C[36] );


HalfAdder fif3fa1( Fou4_S[1], Fou4_C[0], Fif3_S[0], Fif3_C[0] );
FullAdder fif3fa2( Fou4_S[2], Fou4_C[1], pp18[0], Fif3_S[1], Fif3_C[1] );
FullAdder fif3fa3( Fou4_S[3], Fou4_C[2], Fir7_S_[0], Fif3_S[2], Fif3_C[2] );
FullAdder fif3fa4( Fou4_S[4], Fou4_C[3], Sec7_S[0], Fif3_S[3], Fif3_C[3] );
FullAdder fif3fa5( Fou4_S[5], Fou4_C[4], Thi5_S_[0], Fif3_S[4], Fif3_C[4] );
FullAdder fif3fa6( Fou4_S[6], Fou4_C[5], Fou5_S[0], Fif3_S[5], Fif3_C[5] );
FullAdder fif3fa7( Fou4_S[7], Fou4_C[6], Fou5_S[1], Fif3_S[6], Fif3_C[6] );
FullAdder fif3fa8( Fou4_S[8], Fou4_C[7], Fou5_S[2], Fif3_S[7], Fif3_C[7] );
FullAdder fif3fa9( Fou4_S[9], Fou4_C[8], Fou5_S[3], Fif3_S[8], Fif3_C[8] );
FullAdder fif3fa10( Fou4_S[10], Fou4_C[9], Fou5_S[4], Fif3_S[9], Fif3_C[9] );
FullAdder fif3fa11( Fou4_S[11], Fou4_C[10], Fou5_S[5], Fif3_S[10], Fif3_C[10] );
FullAdder fif3fa12( Fou4_S[12], Fou4_C[11], Fou5_S[6], Fif3_S[11], Fif3_C[11] );
FullAdder fif3fa13( Fou4_S[13], Fou4_C[12], Fou5_S[7], Fif3_S[12], Fif3_C[12] );
FullAdder fif3fa14( Fou4_S[14], Fou4_C[13], Fou5_S[8], Fif3_S[13], Fif3_C[13] );
FullAdder fif3fa15( Fou4_S[15], Fou4_C[14], Fou5_S[9], Fif3_S[14], Fif3_C[14] );
FullAdder fif3fa16( Fou4_S[16], Fou4_C[15], Fou5_S[10], Fif3_S[15], Fif3_C[15] );
FullAdder fif3fa17( Fou4_S[17], Fou4_C[16], Fou5_S[11], Fif3_S[16], Fif3_C[16] );
FullAdder fif3fa18( Fou4_S[18], Fou4_C[17], Fou5_S[12], Fif3_S[17], Fif3_C[17] );
FullAdder fif3fa19( Fou4_S[19], Fou4_C[18], Fou5_S[13], Fif3_S[18], Fif3_C[18] );
FullAdder fif3fa20( Fou4_S[20], Fou4_C[19], Fou5_S[14], Fif3_S[19], Fif3_C[19] );
FullAdder fif3fa21( Fou4_S[21], Fou4_C[20], Fou5_S[15], Fif3_S[20], Fif3_C[20] );
FullAdder fif3fa22( Fou4_S[22], Fou4_C[21], Fou5_S[16], Fif3_S[21], Fif3_C[21] );
FullAdder fif3fa23( Fou4_S[23], Fou4_C[22], Fou5_S[17], Fif3_S[22], Fif3_C[22] );
FullAdder fif3fa24( Fou4_S[24], Fou4_C[23], Fou5_S[18], Fif3_S[23], Fif3_C[23] );
FullAdder fif3fa25( Fou4_S[25], Fou4_C[24], Fou5_S[19], Fif3_S[24], Fif3_C[24] );
FullAdder fif3fa26( Fou4_S[26], Fou4_C[25], Fou5_S[20], Fif3_S[25], Fif3_C[25] );
FullAdder fif3fa27( Fou4_S[27], Fou4_C[26], Fou5_S[21], Fif3_S[26], Fif3_C[26] );
FullAdder fif3fa28( Fou4_S[28], Fou4_C[27], Fou5_S[22], Fif3_S[27], Fif3_C[27] );
FullAdder fif3fa29( Fou4_S[29], Fou4_C[28], Fou5_S[23], Fif3_S[28], Fif3_C[28] );
FullAdder fif3fa30( Fou4_S[30], Fou4_C[29], Fou5_S[24], Fif3_S[29], Fif3_C[29] );
FullAdder fif3fa31( Fou4_S[31], Fou4_C[30], Fou5_S[25], Fif3_S[30], Fif3_C[30] );
FullAdder fif3fa32( Fou4_S[32], Fou4_C[31], Fou5_S[26], Fif3_S[31], Fif3_C[31] );
FullAdder fif3fa33( Fou4_S[33], Fou4_C[32], Fou5_S[27], Fif3_S[32], Fif3_C[32] );
HalfAdder fif3fa34( Fou4_C[33], Fou5_S[28], Fif3_S[33], Fif3_C[33] );


HalfAdder fif4fa1( Thi6_S_[0], Fou5_C[1], Fif4_S[0], Fif4_C[0] );
HalfAdder fif4fa2( Fou6_S[0], Fou5_C[2], Fif4_S[1], Fif4_C[1] );
FullAdder fif4fa3( Fou6_S[1], Fou5_C[3], Fou6_C[0], Fif4_S[2], Fif4_C[2] );
FullAdder fif4fa4( Fou6_S[2], Fou5_C[4], Fou6_C[1], Fif4_S[3], Fif4_C[3] );
FullAdder fif4fa5( Fou6_S[3], Fou5_C[5], Fou6_C[2], Fif4_S[4], Fif4_C[4] );
FullAdder fif4fa6( Fou6_S[4], Fou5_C[6], Fou6_C[3], Fif4_S[5], Fif4_C[5] );
FullAdder fif4fa7( Fou6_S[5], Fou5_C[7], Fou6_C[4], Fif4_S[6], Fif4_C[6] );
FullAdder fif4fa8( Fou6_S[6], Fou5_C[8], Fou6_C[5], Fif4_S[7], Fif4_C[7] );
FullAdder fif4fa9( Fou6_S[7], Fou5_C[9], Fou6_C[6], Fif4_S[8], Fif4_C[8] );
FullAdder fif4fa10( Fou6_S[8], Fou5_C[10], Fou6_C[7], Fif4_S[9], Fif4_C[9] );
FullAdder fif4fa11( Fou6_S[9], Fou5_C[11], Fou6_C[8], Fif4_S[10], Fif4_C[10] );
FullAdder fif4fa12( Fou6_S[10], Fou5_C[12], Fou6_C[9], Fif4_S[11], Fif4_C[11] );
FullAdder fif4fa13( Fou6_S[11], Fou5_C[13], Fou6_C[10], Fif4_S[12], Fif4_C[12] );
FullAdder fif4fa14( Fou6_S[12], Fou5_C[14], Fou6_C[11], Fif4_S[13], Fif4_C[13] );
FullAdder fif4fa15( Fou6_S[13], Fou5_C[15], Fou6_C[12], Fif4_S[14], Fif4_C[14] );
FullAdder fif4fa16( Fou6_S[14], Fou5_C[16], Fou6_C[13], Fif4_S[15], Fif4_C[15] );
FullAdder fif4fa17( Fou6_S[15], Fou5_C[17], Fou6_C[14], Fif4_S[16], Fif4_C[16] );
FullAdder fif4fa18( Fou6_S[16], Fou5_C[18], Fou6_C[15], Fif4_S[17], Fif4_C[17] );
FullAdder fif4fa19( Fou6_S[17], Fou5_C[19], Fou6_C[16], Fif4_S[18], Fif4_C[18] );
FullAdder fif4fa20( Fou6_S[18], Fou5_C[20], Fou6_C[17], Fif4_S[19], Fif4_C[19] );
FullAdder fif4fa21( Fou6_S[19], Fou5_C[21], Fou6_C[18], Fif4_S[20], Fif4_C[20] );
FullAdder fif4fa22( Fou6_S[20], Fou5_C[22], Fou6_C[19], Fif4_S[21], Fif4_C[21] );
FullAdder fif4fa23( Fou6_S[21], Fou5_C[23], Fou6_C[20], Fif4_S[22], Fif4_C[22] );
FullAdder fif4fa24( Fou6_S[22], Fou5_C[24], Fou6_C[21], Fif4_S[23], Fif4_C[23] );
FullAdder fif4fa25( Fou6_S[23], Fou5_C[25], Fou6_C[22], Fif4_S[24], Fif4_C[24] );
FullAdder fif4fa26( Fou6_S[24], Fou5_C[26], Fou6_C[23], Fif4_S[25], Fif4_C[25] );
FullAdder fif4fa27( Fou6_S[25], Fou5_C[27], Fou6_C[24], Fif4_S[26], Fif4_C[26] );
FullAdder fif4fa28( Fou6_S[26], Fou5_C[28], Fou6_C[25], Fif4_S[27], Fif4_C[27] );
FullAdder fif4fa29( Fou6_S[27], Fou5_C[29], Fou6_C[26], Fif4_S[28], Fif4_C[28] );
FullAdder fif4fa30( Fou6_S[28], Fou5_C[30], Fou6_C[27], Fif4_S[29], Fif4_C[29] );
FullAdder fif4fa31( Fou6_S[29], Fou5_C[31], Fou6_C[28], Fif4_S[30], Fif4_C[30] );
HalfAdder fif4fa32( Fou6_S[30], Fou6_C[29], Fif4_S[31], Fif4_C[31] );
HalfAdder fif4fa33( Fou6_S[31], Fou6_C[30], Fif4_S[32], Fif4_C[32] );
HalfAdder fif4fa34( Fou6_S[32], Fou6_C[31], Fif4_S[33], Fif4_C[33] );
HalfAdder fif4fa35( Fou6_S[33], Fou6_C[32], Fif4_S[34], Fif4_C[34] );


HalfAdder fif5fa1( Fou7_S[1], Fou7_C[0], Fif5_S[0], Fif5_C[0] );
FullAdder fif5fa2( Fou7_S[2], Fou7_C[1], Sec11_C[0], Fif5_S[1], Fif5_C[1] );
FullAdder fif5fa3( Fou7_S[3], Fou7_C[2], Sec11_C[1], Fif5_S[2], Fif5_C[2] );
FullAdder fif5fa4( Fou7_S[4], Fou7_C[3], Sec11_C[2], Fif5_S[3], Fif5_C[3] );
FullAdder fif5fa5( Fou7_S[5], Fou7_C[4], Sec11_C[3], Fif5_S[4], Fif5_C[4] );
FullAdder fif5fa6( Fou7_S[6], Fou7_C[5], Sec11_C[4], Fif5_S[5], Fif5_C[5] );
FullAdder fif5fa7( Fou7_S[7], Fou7_C[6], Sec11_C[5], Fif5_S[6], Fif5_C[6] );
FullAdder fif5fa8( Fou7_S[8], Fou7_C[7], Sec11_C[6], Fif5_S[7], Fif5_C[7] );
FullAdder fif5fa9( Fou7_S[9], Fou7_C[8], Sec11_C[7], Fif5_S[8], Fif5_C[8] );
FullAdder fif5fa10( Fou7_S[10], Fou7_C[9], Sec11_C[8], Fif5_S[9], Fif5_C[9] );
FullAdder fif5fa11( Fou7_S[11], Fou7_C[10], Sec11_C[9], Fif5_S[10], Fif5_C[10] );
FullAdder fif5fa12( Fou7_S[12], Fou7_C[11], Sec11_C[10], Fif5_S[11], Fif5_C[11] );
FullAdder fif5fa13( Fou7_S[13], Fou7_C[12], Sec11_C[11], Fif5_S[12], Fif5_C[12] );
FullAdder fif5fa14( Fou7_S[14], Fou7_C[13], Sec11_C[12], Fif5_S[13], Fif5_C[13] );
FullAdder fif5fa15( Fou7_S[15], Fou7_C[14], Sec11_C[13], Fif5_S[14], Fif5_C[14] );
FullAdder fif5fa16( Fou7_S[16], Fou7_C[15], Sec11_C[14], Fif5_S[15], Fif5_C[15] );
FullAdder fif5fa17( Fou7_S[17], Fou7_C[16], Sec11_C[15], Fif5_S[16], Fif5_C[16] );
FullAdder fif5fa18( Fou7_S[18], Fou7_C[17], Sec11_C[16], Fif5_S[17], Fif5_C[17] );
FullAdder fif5fa19( Fou7_S[19], Fou7_C[18], Sec11_C[17], Fif5_S[18], Fif5_C[18] );
FullAdder fif5fa20( Fou7_S[20], Fou7_C[19], Sec11_C[18], Fif5_S[19], Fif5_C[19] );
FullAdder fif5fa21( Fou7_S[21], Fou7_C[20], Sec11_C[19], Fif5_S[20], Fif5_C[20] );
FullAdder fif5fa22( Fou7_S[22], Fou7_C[21], Sec11_C[20], Fif5_S[21], Fif5_C[21] );
FullAdder fif5fa23( Fou7_S[23], Fou7_C[22], Sec11_C[21], Fif5_S[22], Fif5_C[22] );
FullAdder fif5fa24( Fou7_S[24], Fou7_C[23], Sec11_C[22], Fif5_S[23], Fif5_C[23] );
FullAdder fif5fa25( Fou7_S[25], Fou7_C[24], Sec11_C[23], Fif5_S[24], Fif5_C[24] );
FullAdder fif5fa26( Fou7_S[26], Fou7_C[25], Sec11_C[24], Fif5_S[25], Fif5_C[25] );
FullAdder fif5fa27( Fou7_S[27], Fou7_C[26], Sec11_C[25], Fif5_S[26], Fif5_C[26] );
FullAdder fif5fa28( Fou7_S[28], Fou7_C[27], Sec11_C[26], Fif5_S[27], Fif5_C[27] );
FullAdder fif5fa29( Fou7_S[29], Fou7_C[28], Sec11_C[27], Fif5_S[28], Fif5_C[28] );
FullAdder fif5fa30( Fou7_S[30], Fou7_C[29], Sec11_C[28], Fif5_S[29], Fif5_C[29] );
FullAdder fif5fa31( Fou7_S[31], Fou7_C[30], Sec11_C[29], Fif5_S[30], Fif5_C[30] );
HalfAdder fif5fa32( Fou7_C[31], Sec11_C[30], Fif5_S[31], Fif5_C[31] );


reg	[31: 0]	Fif1_S_, Fif1_C_;
reg	[36: 0]	Fif2_S_, Fif2_C_;
reg	[33: 0]	Fif3_S_, Fif3_C_;
reg	[34: 0]	Fif4_S_, Fif4_C_;
reg	[31: 0]	Fif5_S_, Fif5_C_;


reg done4;
reg state_done4;

always @(posedge clk or posedge reset) begin
    if (reset) begin
        Fif1_S_ <= 32'b0; Fif1_C_ <= 32'b0;
        Fif2_S_ <= 37'b0; Fif2_C_ <= 37'b0;
        Fif3_S_ <= 34'b0; Fif3_C_ <= 34'b0;
        Fif4_S_ <= 35'b0; Fif4_C_ <= 35'b0;
        Fif5_S_ <= 32'b0; Fif5_C_ <= 32'b0;
        done4   <= 1'b0;
        state_done4 <= 1'b0;
    end else begin
        case (state_done4)
            1'b0: begin
                if (done3) begin
                    Fif1_S_ <= Fif1_S; Fif1_C_ <= Fif1_C;
                    Fif2_S_ <= Fif2_S; Fif2_C_ <= Fif2_C;
                    Fif3_S_ <= Fif3_S; Fif3_C_ <= Fif3_C;
                    Fif4_S_ <= Fif4_S; Fif4_C_ <= Fif4_C;
                    Fif5_S_ <= Fif5_S; Fif5_C_ <= Fif5_C;
                    done4 <= 1'b1;
                    state_done4 <= 1'b1;
                end else begin
                    done4 <= 1'b0;
                end
            end
            1'b1: begin
                done4 <= 1'b0;
                if (!done3)
                    state_done4 <= 1'b0;
            end
        endcase
    end
end


//===================Sixth stage===============================


wire	[31: 0]	Six1_S_, Six1_C_;
wire	[35: 0]	Six2_S_, Six2_C_;
wire	[33: 0]	Six3_S_, Six3_C_;
wire	[34: 0]	Six4_S_, Six4_C_;
wire	[31: 0]	Six5_S_, Six5_C_;


assign Six1_S_ = Fif1_S_;
assign Six1_C_ = Fif1_C_;


HalfAdder six2fa1( Fif2_S_[1], Fif2_C_[0], Six2_S_[0], Six2_C_[0] );
HalfAdder six2fa2( Fif2_S_[2], Fif2_C_[1], Six2_S_[1], Six2_C_[1] );
HalfAdder six2fa3( Fif2_S_[3], Fif2_C_[2], Six2_S_[2], Six2_C_[2] );
HalfAdder six2fa4( Fif2_S_[4], Fif2_C_[3], Six2_S_[3], Six2_C_[3] );
HalfAdder six2fa5( Fif2_S_[5], Fif2_C_[4], Six2_S_[4], Six2_C_[4] );
HalfAdder six2fa6( Fif2_S_[6], Fif2_C_[5], Six2_S_[5], Six2_C_[5] );
HalfAdder six2fa7( Fif2_S_[7], Fif2_C_[6], Six2_S_[6], Six2_C_[6] );
HalfAdder six2fa8( Fif2_S_[8], Fif2_C_[7], Six2_S_[7], Six2_C_[7] );
HalfAdder six2fa9( Fif2_S_[9], Fif2_C_[8], Six2_S_[8], Six2_C_[8] );
HalfAdder six2fa10( Fif2_S_[10], Fif2_C_[9], Six2_S_[9], Six2_C_[9] );
HalfAdder six2fa11( Fif2_S_[11], Fif2_C_[10], Six2_S_[10], Six2_C_[10] );
HalfAdder six2fa12( Fif2_S_[12], Fif2_C_[11], Six2_S_[11], Six2_C_[11] );
HalfAdder six2fa13( Fif2_S_[13], Fif2_C_[12], Six2_S_[12], Six2_C_[12] );
HalfAdder six2fa14( Fif2_S_[14], Fif2_C_[13], Six2_S_[13], Six2_C_[13] );
HalfAdder six2fa15( Fif2_S_[15], Fif2_C_[14], Six2_S_[14], Six2_C_[14] );
HalfAdder six2fa16( Fif2_S_[16], Fif2_C_[15], Six2_S_[15], Six2_C_[15] );
HalfAdder six2fa17( Fif2_S_[17], Fif2_C_[16], Six2_S_[16], Six2_C_[16] );
HalfAdder six2fa18( Fif2_S_[18], Fif2_C_[17], Six2_S_[17], Six2_C_[17] );
HalfAdder six2fa19( Fif2_S_[19], Fif2_C_[18], Six2_S_[18], Six2_C_[18] );
HalfAdder six2fa20( Fif2_S_[20], Fif2_C_[19], Six2_S_[19], Six2_C_[19] );
HalfAdder six2fa21( Fif2_S_[21], Fif2_C_[20], Six2_S_[20], Six2_C_[20] );
HalfAdder six2fa22( Fif2_S_[22], Fif2_C_[21], Six2_S_[21], Six2_C_[21] );
HalfAdder six2fa23( Fif2_S_[23], Fif2_C_[22], Six2_S_[22], Six2_C_[22] );
HalfAdder six2fa24( Fif2_S_[24], Fif2_C_[23], Six2_S_[23], Six2_C_[23] );
HalfAdder six2fa25( Fif2_S_[25], Fif2_C_[24], Six2_S_[24], Six2_C_[24] );
HalfAdder six2fa26( Fif2_S_[26], Fif2_C_[25], Six2_S_[25], Six2_C_[25] );
HalfAdder six2fa27( Fif2_S_[27], Fif2_C_[26], Six2_S_[26], Six2_C_[26] );
FullAdder six2fa28( Fou2_S[30], Fif2_S_[28], Fif2_C_[27], Six2_S_[27], Six2_C_[27] );
FullAdder six2fa29( Fou2_S[31], Fif2_S_[29], Fif2_C_[28], Six2_S_[28], Six2_C_[28] );
FullAdder six2fa30( Fou2_S[32], Fif2_S_[30], Fif2_C_[29], Six2_S_[29], Six2_C_[29] );
FullAdder six2fa31( Fou2_S[33], Fif2_S_[31], Fif2_C_[30], Six2_S_[30], Six2_C_[30] );
HalfAdder six2fa32( Fif2_S_[32], Fif2_C_[31], Six2_S_[31], Six2_C_[31] );
HalfAdder six2fa33( Fif2_S_[33], Fif2_C_[32], Six2_S_[32], Six2_C_[32] );
HalfAdder six2fa34( Fif2_S_[34], Fif2_C_[33], Six2_S_[33], Six2_C_[33] );
HalfAdder six2fa35( Fif2_S_[35], Fif2_C_[34], Six2_S_[34], Six2_C_[34] );
HalfAdder six2fa36( Fif2_S_[36], Fif2_C_[35], Six2_S_[35], Six2_C_[35] );

assign Six3_S_ = Fif3_S_;
assign Six3_C_ = Fif3_C_;


HalfAdder six4fa1( Fif4_S_[1], Fif4_C_[0], Six4_S_[0], Six4_C_[0] );
HalfAdder six4fa2( Fif4_S_[2], Fif4_C_[1], Six4_S_[1], Six4_C_[1] );
HalfAdder six4fa3( Fif4_S_[3], Fif4_C_[2], Six4_S_[2], Six4_C_[2] );
HalfAdder six4fa4( Fif4_S_[4], Fif4_C_[3], Six4_S_[3], Six4_C_[3] );
HalfAdder six4fa5( Fif4_S_[5], Fif4_C_[4], Six4_S_[4], Six4_C_[4] );
HalfAdder six4fa6( Fif4_S_[6], Fif4_C_[5], Six4_S_[5], Six4_C_[5] );
HalfAdder six4fa7( Fif4_S_[7], Fif4_C_[6], Six4_S_[6], Six4_C_[6] );
HalfAdder six4fa8( Fif4_S_[8], Fif4_C_[7], Six4_S_[7], Six4_C_[7] );
HalfAdder six4fa9( Fif4_S_[9], Fif4_C_[8], Six4_S_[8], Six4_C_[8] );
HalfAdder six4fa10( Fif4_S_[10], Fif4_C_[9], Six4_S_[9], Six4_C_[9] );
HalfAdder six4fa11( Fif4_S_[11], Fif4_C_[10], Six4_S_[10], Six4_C_[10] );
HalfAdder six4fa12( Fif4_S_[12], Fif4_C_[11], Six4_S_[11], Six4_C_[11] );
HalfAdder six4fa13( Fif4_S_[13], Fif4_C_[12], Six4_S_[12], Six4_C_[12] );
HalfAdder six4fa14( Fif4_S_[14], Fif4_C_[13], Six4_S_[13], Six4_C_[13] );
HalfAdder six4fa15( Fif4_S_[15], Fif4_C_[14], Six4_S_[14], Six4_C_[14] );
HalfAdder six4fa16( Fif4_S_[16], Fif4_C_[15], Six4_S_[15], Six4_C_[15] );
HalfAdder six4fa17( Fif4_S_[17], Fif4_C_[16], Six4_S_[16], Six4_C_[16] );
HalfAdder six4fa18( Fif4_S_[18], Fif4_C_[17], Six4_S_[17], Six4_C_[17] );
HalfAdder six4fa19( Fif4_S_[19], Fif4_C_[18], Six4_S_[18], Six4_C_[18] );
HalfAdder six4fa20( Fif4_S_[20], Fif4_C_[19], Six4_S_[19], Six4_C_[19] );
HalfAdder six4fa21( Fif4_S_[21], Fif4_C_[20], Six4_S_[20], Six4_C_[20] );
HalfAdder six4fa22( Fif4_S_[22], Fif4_C_[21], Six4_S_[21], Six4_C_[21] );
HalfAdder six4fa23( Fif4_S_[23], Fif4_C_[22], Six4_S_[22], Six4_C_[22] );
HalfAdder six4fa24( Fif4_S_[24], Fif4_C_[23], Six4_S_[23], Six4_C_[23] );
HalfAdder six4fa25( Fif4_S_[25], Fif4_C_[24], Six4_S_[24], Six4_C_[24] );
HalfAdder six4fa26( Fif4_S_[26], Fif4_C_[25], Six4_S_[25], Six4_C_[25] );
FullAdder six4fa27( Fou5_S[29], Fif4_S_[27], Fif4_C_[26], Six4_S_[26], Six4_C_[26] );
FullAdder six4fa28( Fou5_S[30], Fif4_S_[28], Fif4_C_[27], Six4_S_[27], Six4_C_[27] );
FullAdder six4fa29( Fou5_S[31], Fif4_S_[29], Fif4_C_[28], Six4_S_[28], Six4_C_[28] );
FullAdder six4fa30( Sec8_S[31], Fif4_S_[30], Fif4_C_[29], Six4_S_[29], Six4_C_[29] );
HalfAdder six4fa31( Fif4_S_[31], Fif4_C_[30], Six4_S_[30], Six4_C_[30] );
HalfAdder six4fa32( Fif4_S_[32], Fif4_C_[31], Six4_S_[31], Six4_C_[31] );
HalfAdder six4fa33( Fif4_S_[33], Fif4_C_[32], Six4_S_[32], Six4_C_[32] );
HalfAdder six4fa34( Fif4_S_[34], Fif4_C_[33], Six4_S_[33], Six4_C_[33] );
HalfAdder six4fa35( Fou6_C[33], Fif4_C_[34], Six4_S_[34], Six4_C_[34] );


assign Six5_S_ = Fif5_S_;
assign Six5_C_ = Fif5_C_;


reg	[31: 0]	Six1_S, Six1_C;
reg	[35: 0]	Six2_S, Six2_C;
reg	[33: 0]	Six3_S, Six3_C;
reg	[34: 0]	Six4_S, Six4_C;
reg	[31: 0]	Six5_S, Six5_C;


reg done5;
reg state_done5;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Six1_S <= 32'b0;  Six1_C <= 32'b0;
    Six2_S <= 36'b0;  Six2_C <= 36'b0;
    Six3_S <= 34'b0;  Six3_C <= 34'b0;
    Six4_S <= 35'b0;  Six4_C <= 35'b0;
    Six5_S <= 32'b0;  Six5_C <= 32'b0;
    done5 <= 1'b0;
    state_done5 <= 1'b0;
  end else begin
    case (state_done5)
      1'b0: begin
        if (done4) begin
          Six1_S <= Six1_S_;  Six1_C <= Six1_C_;
          Six2_S <= Six2_S_;  Six2_C <= Six2_C_;
          Six3_S <= Six3_S_;  Six3_C <= Six3_C_;
          Six4_S <= Six4_S_;  Six4_C <= Six4_C_;
          Six5_S <= Six5_S_;  Six5_C <= Six5_C_;
          done5 <= 1'b1;
          state_done5 <= 1'b1;
        end else begin
          done5 <= 1'b0;
        end
      end
      1'b1: begin
        done5 <= 1'b0;
        if (!done4)
          state_done5 <= 1'b0;
      end
    endcase
  end
end


//===================Seventh stage===============================


wire	[31: 0]	Sev1_S, Sev1_C;
wire	[35: 0]	Sev2_S, Sev2_C;
wire	[34: 0]	Sev3_S, Sev3_C;

HalfAdder sev1fa1( Six1_S[1], Six1_C[0], Sev1_S[0], Sev1_C[0] );
HalfAdder sev1fa2( Six1_S[2], Six1_C[1], Sev1_S[1], Sev1_C[1] );
FullAdder sev1fa3( Fou2_C[0], Six1_S[3], Six1_C[2], Sev1_S[2], Sev1_C[2] );
FullAdder sev1fa4( Fif2_S_[0], Six1_S[4], Six1_C[3], Sev1_S[3], Sev1_C[3] );
FullAdder sev1fa5( Six2_S[0], Six1_S[5], Six1_C[4], Sev1_S[4], Sev1_C[4] );
FullAdder sev1fa6( Six2_S[1], Six1_S[6], Six1_C[5], Sev1_S[5], Sev1_C[5] );
FullAdder sev1fa7( Six2_S[2], Six1_S[7], Six1_C[6], Sev1_S[6], Sev1_C[6] );
FullAdder sev1fa8( Six2_S[3], Six1_S[8], Six1_C[7], Sev1_S[7], Sev1_C[7] );
FullAdder sev1fa9( Six2_S[4], Six1_S[9], Six1_C[8], Sev1_S[8], Sev1_C[8] );
FullAdder sev1fa10( Six2_S[5], Six1_S[10], Six1_C[9], Sev1_S[9], Sev1_C[9] );
FullAdder sev1fa11( Six2_S[6], Six1_S[11], Six1_C[10], Sev1_S[10], Sev1_C[10] );
FullAdder sev1fa12( Six2_S[7], Six1_S[12], Six1_C[11], Sev1_S[11], Sev1_C[11] );
FullAdder sev1fa13( Six2_S[8], Six1_S[13], Six1_C[12], Sev1_S[12], Sev1_C[12] );
FullAdder sev1fa14( Six2_S[9], Six1_S[14], Six1_C[13], Sev1_S[13], Sev1_C[13] );
FullAdder sev1fa15( Six2_S[10], Six1_S[15], Six1_C[14], Sev1_S[14], Sev1_C[14] );
FullAdder sev1fa16( Six2_S[11], Six1_S[16], Six1_C[15], Sev1_S[15], Sev1_C[15] );
FullAdder sev1fa17( Six2_S[12], Six1_S[17], Six1_C[16], Sev1_S[16], Sev1_C[16] );
FullAdder sev1fa18( Six2_S[13], Six1_S[18], Six1_C[17], Sev1_S[17], Sev1_C[17] );
FullAdder sev1fa19( Six2_S[14], Six1_S[19], Six1_C[18], Sev1_S[18], Sev1_C[18] );
FullAdder sev1fa20( Six2_S[15], Six1_S[20], Six1_C[19], Sev1_S[19], Sev1_C[19] );
FullAdder sev1fa21( Six2_S[16], Six1_S[21], Six1_C[20], Sev1_S[20], Sev1_C[20] );
FullAdder sev1fa22( Six2_S[17], Six1_S[22], Six1_C[21], Sev1_S[21], Sev1_C[21] );
FullAdder sev1fa23( Six2_S[18], Six1_S[23], Six1_C[22], Sev1_S[22], Sev1_C[22] );
FullAdder sev1fa24( Six2_S[19], Six1_S[24], Six1_C[23], Sev1_S[23], Sev1_C[23] );
FullAdder sev1fa25( Six2_S[20], Six1_S[25], Six1_C[24], Sev1_S[24], Sev1_C[24] );
FullAdder sev1fa26( Six2_S[21], Six1_S[26], Six1_C[25], Sev1_S[25], Sev1_C[25] );
FullAdder sev1fa27( Six2_S[22], Six1_S[27], Six1_C[26], Sev1_S[26], Sev1_C[26] );
FullAdder sev1fa28( Six2_S[23], Six1_S[28], Six1_C[27], Sev1_S[27], Sev1_C[27] );
FullAdder sev1fa29( Six2_S[24], Six1_S[29], Six1_C[28], Sev1_S[28], Sev1_C[28] );
FullAdder sev1fa30( Six2_S[25], Six1_S[30], Six1_C[29], Sev1_S[29], Sev1_C[29] );
FullAdder sev1fa31( Six2_S[26], Six1_S[31], Six1_C[30], Sev1_S[30], Sev1_C[30] );
HalfAdder sev1fa32( Six2_S[27], Six1_C[31], Sev1_S[31], Sev1_C[31] );



HalfAdder sev2fa1( Thi4_S_[0], Six2_C[4], Sev2_S[0], Sev2_C[0] );
HalfAdder sev2fa2( Fou4_S[0], Six2_C[5], Sev2_S[1], Sev2_C[1] );
HalfAdder sev2fa3( Six3_S[0], Six2_C[6], Sev2_S[2], Sev2_C[2] );
FullAdder sev2fa4( Six3_S[1], Six2_C[7], Six3_C[0], Sev2_S[3], Sev2_C[3] );
FullAdder sev2fa5( Six3_S[2], Six2_C[8], Six3_C[1], Sev2_S[4], Sev2_C[4] );
FullAdder sev2fa6( Six3_S[3], Six2_C[9], Six3_C[2], Sev2_S[5], Sev2_C[5] );
FullAdder sev2fa7( Six3_S[4], Six2_C[10], Six3_C[3], Sev2_S[6], Sev2_C[6] );
FullAdder sev2fa8( Six3_S[5], Six2_C[11], Six3_C[4], Sev2_S[7], Sev2_C[7] );
FullAdder sev2fa9( Six3_S[6], Six2_C[12], Six3_C[5], Sev2_S[8], Sev2_C[8] );
FullAdder sev2fa10( Six3_S[7], Six2_C[13], Six3_C[6], Sev2_S[9], Sev2_C[9] );
FullAdder sev2fa11( Six3_S[8], Six2_C[14], Six3_C[7], Sev2_S[10], Sev2_C[10] );
FullAdder sev2fa12( Six3_S[9], Six2_C[15], Six3_C[8], Sev2_S[11], Sev2_C[11] );
FullAdder sev2fa13( Six3_S[10], Six2_C[16], Six3_C[9], Sev2_S[12], Sev2_C[12] );
FullAdder sev2fa14( Six3_S[11], Six2_C[17], Six3_C[10], Sev2_S[13], Sev2_C[13] );
FullAdder sev2fa15( Six3_S[12], Six2_C[18], Six3_C[11], Sev2_S[14], Sev2_C[14] );
FullAdder sev2fa16( Six3_S[13], Six2_C[19], Six3_C[12], Sev2_S[15], Sev2_C[15] );
FullAdder sev2fa17( Six3_S[14], Six2_C[20], Six3_C[13], Sev2_S[16], Sev2_C[16] );
FullAdder sev2fa18( Six3_S[15], Six2_C[21], Six3_C[14], Sev2_S[17], Sev2_C[17] );
FullAdder sev2fa19( Six3_S[16], Six2_C[22], Six3_C[15], Sev2_S[18], Sev2_C[18] );
FullAdder sev2fa20( Six3_S[17], Six2_C[23], Six3_C[16], Sev2_S[19], Sev2_C[19] );
FullAdder sev2fa21( Six3_S[18], Six2_C[24], Six3_C[17], Sev2_S[20], Sev2_C[20] );
FullAdder sev2fa22( Six3_S[19], Six2_C[25], Six3_C[18], Sev2_S[21], Sev2_C[21] );
FullAdder sev2fa23( Six3_S[20], Six2_C[26], Six3_C[19], Sev2_S[22], Sev2_C[22] );
FullAdder sev2fa24( Six3_S[21], Six2_C[27], Six3_C[20], Sev2_S[23], Sev2_C[23] );
FullAdder sev2fa25( Six3_S[22], Six2_C[28], Six3_C[21], Sev2_S[24], Sev2_C[24] );
FullAdder sev2fa26( Six3_S[23], Six2_C[29], Six3_C[22], Sev2_S[25], Sev2_C[25] );
FullAdder sev2fa27( Six3_S[24], Six2_C[30], Six3_C[23], Sev2_S[26], Sev2_C[26] );
FullAdder sev2fa28( Six3_S[25], Six2_C[31], Six3_C[24], Sev2_S[27], Sev2_C[27] );
FullAdder sev2fa29( Six3_S[26], Six2_C[32], Six3_C[25], Sev2_S[28], Sev2_C[28] );
FullAdder sev2fa30( Six3_S[27], Six2_C[33], Six3_C[26], Sev2_S[29], Sev2_C[29] );
FullAdder sev2fa31( Six3_S[28], Six2_C[34], Six3_C[27], Sev2_S[30], Sev2_C[30] );
FullAdder sev2fa32( Six3_S[29], Six2_C[35], Six3_C[28], Sev2_S[31], Sev2_C[31] );
HalfAdder sev2fa33( Six3_S[30], Six3_C[29], Sev2_S[32], Sev2_C[32] );
HalfAdder sev2fa34( Six3_S[31], Six3_C[30], Sev2_S[33], Sev2_C[33] );
HalfAdder sev2fa35( Six3_S[32], Six3_C[31], Sev2_S[34], Sev2_C[34] );
HalfAdder sev2fa36( Six3_S[33], Six3_C[32], Sev2_S[35], Sev2_C[35] );

HalfAdder sev3fa1( Six4_S[1], Six4_C[0], Sev3_S[0], Sev3_C[0] );
FullAdder sev3fa2( Six4_S[2], Six4_C[1], pp27[0], Sev3_S[1], Sev3_C[1] );
FullAdder sev3fa3( Six4_S[3], Six4_C[2], Fir10_S_[0], Sev3_S[2], Sev3_C[2] );
FullAdder sev3fa4( Six4_S[4], Six4_C[3], Sec10_S[0], Sev3_S[3], Sev3_C[3] );
FullAdder sev3fa5( Six4_S[5], Six4_C[4], Thi7_S_[0], Sev3_S[4], Sev3_C[4] );
FullAdder sev3fa6( Six4_S[6], Six4_C[5], Fou7_S[0], Sev3_S[5], Sev3_C[5] );
FullAdder sev3fa7( Six4_S[7], Six4_C[6], Six5_S[0], Sev3_S[6], Sev3_C[6] );
FullAdder sev3fa8( Six4_S[8], Six4_C[7], Six5_S[1], Sev3_S[7], Sev3_C[7] );
FullAdder sev3fa9( Six4_S[9], Six4_C[8], Six5_S[2], Sev3_S[8], Sev3_C[8] );
FullAdder sev3fa10( Six4_S[10], Six4_C[9], Six5_S[3], Sev3_S[9], Sev3_C[9] );
FullAdder sev3fa11( Six4_S[11], Six4_C[10], Six5_S[4], Sev3_S[10], Sev3_C[10] );
FullAdder sev3fa12( Six4_S[12], Six4_C[11], Six5_S[5], Sev3_S[11], Sev3_C[11] );
FullAdder sev3fa13( Six4_S[13], Six4_C[12], Six5_S[6], Sev3_S[12], Sev3_C[12] );
FullAdder sev3fa14( Six4_S[14], Six4_C[13], Six5_S[7], Sev3_S[13], Sev3_C[13] );
FullAdder sev3fa15( Six4_S[15], Six4_C[14], Six5_S[8], Sev3_S[14], Sev3_C[14] );
FullAdder sev3fa16( Six4_S[16], Six4_C[15], Six5_S[9], Sev3_S[15], Sev3_C[15] );
FullAdder sev3fa17( Six4_S[17], Six4_C[16], Six5_S[10], Sev3_S[16], Sev3_C[16] );
FullAdder sev3fa18( Six4_S[18], Six4_C[17], Six5_S[11], Sev3_S[17], Sev3_C[17] );
FullAdder sev3fa19( Six4_S[19], Six4_C[18], Six5_S[12], Sev3_S[18], Sev3_C[18] );
FullAdder sev3fa20( Six4_S[20], Six4_C[19], Six5_S[13], Sev3_S[19], Sev3_C[19] );
FullAdder sev3fa21( Six4_S[21], Six4_C[20], Six5_S[14], Sev3_S[20], Sev3_C[20] );
FullAdder sev3fa22( Six4_S[22], Six4_C[21], Six5_S[15], Sev3_S[21], Sev3_C[21] );
FullAdder sev3fa23( Six4_S[23], Six4_C[22], Six5_S[16], Sev3_S[22], Sev3_C[22] );
FullAdder sev3fa24( Six4_S[24], Six4_C[23], Six5_S[17], Sev3_S[23], Sev3_C[23] );
FullAdder sev3fa25( Six4_S[25], Six4_C[24], Six5_S[18], Sev3_S[24], Sev3_C[24] );
FullAdder sev3fa26( Six4_S[26], Six4_C[25], Six5_S[19], Sev3_S[25], Sev3_C[25] );
FullAdder sev3fa27( Six4_S[27], Six4_C[26], Six5_S[20], Sev3_S[26], Sev3_C[26] );
FullAdder sev3fa28( Six4_S[28], Six4_C[27], Six5_S[21], Sev3_S[27], Sev3_C[27] );
FullAdder sev3fa29( Six4_S[29], Six4_C[28], Six5_S[22], Sev3_S[28], Sev3_C[28] );
FullAdder sev3fa30( Six4_S[30], Six4_C[29], Six5_S[23], Sev3_S[29], Sev3_C[29] );
FullAdder sev3fa31( Six4_S[31], Six4_C[30], Six5_S[24], Sev3_S[30], Sev3_C[30] );
FullAdder sev3fa32( Six4_S[32], Six4_C[31], Six5_S[25], Sev3_S[31], Sev3_C[31] );
FullAdder sev3fa33( Six4_S[33], Six4_C[32], Six5_S[26], Sev3_S[32], Sev3_C[32] );
FullAdder sev3fa34( Six4_S[34], Six4_C[33], Six5_S[27], Sev3_S[33], Sev3_C[33] );
HalfAdder sev3fa35( Six4_C[34], Six5_S[28], Sev3_S[34], Sev3_C[34] );


reg	[31: 0]	Sev1_S_, Sev1_C_;
reg	[35: 0]	Sev2_S_, Sev2_C_;
reg	[34: 0]	Sev3_S_, Sev3_C_;

reg done6;
reg state_done6;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Sev1_S_ <= 32'b0;  Sev1_C_ <= 32'b0;
    Sev2_S_ <= 36'b0;  Sev2_C_ <= 36'b0;
    Sev3_S_ <= 35'b0;  Sev3_C_ <= 35'b0;
    done6 <= 1'b0;
    state_done6 <= 1'b0;
  end else begin
    case (state_done6)
      1'b0: begin
        if (done5) begin
          Sev1_S_ <= Sev1_S;  Sev1_C_ <= Sev1_C;
          Sev2_S_ <= Sev2_S;  Sev2_C_ <= Sev2_C;
          Sev3_S_ <= Sev3_S;  Sev3_C_ <= Sev3_C;
          done6 <= 1'b1;
          state_done6 <= 1'b1;
        end else begin
          done6 <= 1'b0;
        end
      end
      1'b1: begin
        done6 <= 1'b0;
        if (!done5)
          state_done6 <= 1'b0;
      end
    endcase
  end
end


//===================Eighth stage===============================

wire	[31: 0]	Eig1_S_, Eig1_C_;
wire	[35: 0]	Eig2_S_, Eig2_C_;
wire	[36: 0]	Eig3_S_, Eig3_C_;


assign Eig1_S_=Sev1_S_;
assign Eig1_C_=Sev1_C_;

HalfAdder eig2fa1( Sev2_C_[0], Sev2_S_[1], Eig2_S_[0], Eig2_C_[0] );
HalfAdder eig2fa2( Sev2_C_[1], Sev2_S_[2], Eig2_S_[1], Eig2_C_[1] );
HalfAdder eig2fa3( Sev2_C_[2], Sev2_S_[3], Eig2_S_[2], Eig2_C_[2] );
HalfAdder eig2fa4( Sev2_C_[3], Sev2_S_[4], Eig2_S_[3], Eig2_C_[3] );
HalfAdder eig2fa5( Sev2_C_[4], Sev2_S_[5], Eig2_S_[4], Eig2_C_[4] );
HalfAdder eig2fa6( Sev2_C_[5], Sev2_S_[6], Eig2_S_[5], Eig2_C_[5] );
HalfAdder eig2fa7( Sev2_C_[6], Sev2_S_[7], Eig2_S_[6], Eig2_C_[6] );
HalfAdder eig2fa8( Sev2_C_[7], Sev2_S_[8], Eig2_S_[7], Eig2_C_[7] );
HalfAdder eig2fa9( Sev2_C_[8], Sev2_S_[9], Eig2_S_[8], Eig2_C_[8] );
HalfAdder eig2fa10( Sev2_C_[9], Sev2_S_[10], Eig2_S_[9], Eig2_C_[9] );
HalfAdder eig2fa11( Sev2_C_[10], Sev2_S_[11], Eig2_S_[10], Eig2_C_[10] );
HalfAdder eig2fa12( Sev2_C_[11], Sev2_S_[12], Eig2_S_[11], Eig2_C_[11] );
HalfAdder eig2fa13( Sev2_C_[12], Sev2_S_[13], Eig2_S_[12], Eig2_C_[12] );
HalfAdder eig2fa14( Sev2_C_[13], Sev2_S_[14], Eig2_S_[13], Eig2_C_[13] );
HalfAdder eig2fa15( Sev2_C_[14], Sev2_S_[15], Eig2_S_[14], Eig2_C_[14] );
HalfAdder eig2fa16( Sev2_C_[15], Sev2_S_[16], Eig2_S_[15], Eig2_C_[15] );
HalfAdder eig2fa17( Sev2_C_[16], Sev2_S_[17], Eig2_S_[16], Eig2_C_[16] );
HalfAdder eig2fa18( Sev2_C_[17], Sev2_S_[18], Eig2_S_[17], Eig2_C_[17] );
HalfAdder eig2fa19( Sev2_C_[18], Sev2_S_[19], Eig2_S_[18], Eig2_C_[18] );
HalfAdder eig2fa20( Sev2_C_[19], Sev2_S_[20], Eig2_S_[19], Eig2_C_[19] );
HalfAdder eig2fa21( Sev2_C_[20], Sev2_S_[21], Eig2_S_[20], Eig2_C_[20] );
HalfAdder eig2fa22( Sev2_C_[21], Sev2_S_[22], Eig2_S_[21], Eig2_C_[21] );
FullAdder eig2fa23( Six2_S[28], Sev2_C_[22], Sev2_S_[23], Eig2_S_[22], Eig2_C_[22] );
FullAdder eig2fa24( Six2_S[29], Sev2_C_[23], Sev2_S_[24], Eig2_S_[23], Eig2_C_[23] );
FullAdder eig2fa25( Six2_S[30], Sev2_C_[24], Sev2_S_[25], Eig2_S_[24], Eig2_C_[24] );
FullAdder eig2fa26( Six2_S[31], Sev2_C_[25], Sev2_S_[26], Eig2_S_[25], Eig2_C_[25] );
FullAdder eig2fa27( Six2_S[32], Sev2_C_[26], Sev2_S_[27], Eig2_S_[26], Eig2_C_[26] );
FullAdder eig2fa28( Six2_S[33], Sev2_C_[27], Sev2_S_[28], Eig2_S_[27], Eig2_C_[27] );
FullAdder eig2fa29( Six2_S[34], Sev2_C_[28], Sev2_S_[29], Eig2_S_[28], Eig2_C_[28] );
FullAdder eig2fa30( Six2_S[35], Sev2_C_[29], Sev2_S_[30], Eig2_S_[29], Eig2_C_[29] );
FullAdder eig2fa31( Fif2_C_[36], Sev2_C_[30], Sev2_S_[31], Eig2_S_[30], Eig2_C_[30] );
HalfAdder eig2fa32( Sev2_C_[31], Sev2_S_[32], Eig2_S_[31], Eig2_C_[31] );
HalfAdder eig2fa33( Sev2_C_[32], Sev2_S_[33], Eig2_S_[32], Eig2_C_[32] );
HalfAdder eig2fa34( Sev2_C_[33], Sev2_S_[34], Eig2_S_[33], Eig2_C_[33] );
HalfAdder eig2fa35( Sev2_C_[34], Sev2_S_[35], Eig2_S_[34], Eig2_C_[34] );
HalfAdder eig2fa36( Sev2_C_[35], Six3_C[33], Eig2_S_[35], Eig2_C_[35] );

HalfAdder eig3fa1( Sev3_C_[0], Sev3_S_[1], Eig3_S_[0], Eig3_C_[0] );
HalfAdder eig3fa2( Sev3_C_[1], Sev3_S_[2], Eig3_S_[1], Eig3_C_[1] );
HalfAdder eig3fa3( Sev3_C_[2], Sev3_S_[3], Eig3_S_[2], Eig3_C_[2] );
HalfAdder eig3fa4( Sev3_C_[3], Sev3_S_[4], Eig3_S_[3], Eig3_C_[3] );
HalfAdder eig3fa5( Sev3_C_[4], Sev3_S_[5], Eig3_S_[4], Eig3_C_[4] );
HalfAdder eig3fa6( Sev3_C_[5], Sev3_S_[6], Eig3_S_[5], Eig3_C_[5] );
FullAdder eig3fa7( Sev3_C_[6], Sev3_S_[7], Six5_C[0], Eig3_S_[6], Eig3_C_[6] );
FullAdder eig3fa8( Sev3_C_[7], Sev3_S_[8], Six5_C[1], Eig3_S_[7], Eig3_C_[7] );
FullAdder eig3fa9( Sev3_C_[8], Sev3_S_[9], Six5_C[2], Eig3_S_[8], Eig3_C_[8] );
FullAdder eig3fa10( Sev3_C_[9],  Sev3_S_[10], Six5_C[3],  Eig3_S_[9],  Eig3_C_[9] );
FullAdder eig3fa11( Sev3_C_[10], Sev3_S_[11], Six5_C[4],  Eig3_S_[10], Eig3_C_[10] );
FullAdder eig3fa12( Sev3_C_[11], Sev3_S_[12], Six5_C[5],  Eig3_S_[11], Eig3_C_[11] );
FullAdder eig3fa13( Sev3_C_[12], Sev3_S_[13], Six5_C[6],  Eig3_S_[12], Eig3_C_[12] );
FullAdder eig3fa14( Sev3_C_[13], Sev3_S_[14], Six5_C[7],  Eig3_S_[13], Eig3_C_[13] );
FullAdder eig3fa15( Sev3_C_[14], Sev3_S_[15], Six5_C[8],  Eig3_S_[14], Eig3_C_[14] );
FullAdder eig3fa16( Sev3_C_[15], Sev3_S_[16], Six5_C[9],  Eig3_S_[15], Eig3_C_[15] );
FullAdder eig3fa17( Sev3_C_[16], Sev3_S_[17], Six5_C[10], Eig3_S_[16], Eig3_C_[16] );
FullAdder eig3fa18( Sev3_C_[17], Sev3_S_[18], Six5_C[11], Eig3_S_[17], Eig3_C_[17] );
FullAdder eig3fa19( Sev3_C_[18], Sev3_S_[19], Six5_C[12], Eig3_S_[18], Eig3_C_[18] );
FullAdder eig3fa20( Sev3_C_[19], Sev3_S_[20], Six5_C[13], Eig3_S_[19], Eig3_C_[19] );
FullAdder eig3fa21( Sev3_C_[20], Sev3_S_[21], Six5_C[14], Eig3_S_[20], Eig3_C_[20] );
FullAdder eig3fa22( Sev3_C_[21], Sev3_S_[22], Six5_C[15], Eig3_S_[21], Eig3_C_[21] );
FullAdder eig3fa23( Sev3_C_[22], Sev3_S_[23], Six5_C[16], Eig3_S_[22], Eig3_C_[22] );
FullAdder eig3fa24( Sev3_C_[23], Sev3_S_[24], Six5_C[17], Eig3_S_[23], Eig3_C_[23] );
FullAdder eig3fa25( Sev3_C_[24], Sev3_S_[25], Six5_C[18], Eig3_S_[24], Eig3_C_[24] );
FullAdder eig3fa26( Sev3_C_[25], Sev3_S_[26], Six5_C[19], Eig3_S_[25], Eig3_C_[25] );
FullAdder eig3fa27( Sev3_C_[26], Sev3_S_[27], Six5_C[20], Eig3_S_[26], Eig3_C_[26] );
FullAdder eig3fa28( Sev3_C_[27], Sev3_S_[28], Six5_C[21], Eig3_S_[27], Eig3_C_[27] );
FullAdder eig3fa29( Sev3_C_[28], Sev3_S_[29], Six5_C[22], Eig3_S_[28], Eig3_C_[28] );
FullAdder eig3fa30( Sev3_C_[29], Sev3_S_[30], Six5_C[23], Eig3_S_[29], Eig3_C_[29] );
FullAdder eig3fa31( Sev3_C_[30], Sev3_S_[31], Six5_C[24], Eig3_S_[30], Eig3_C_[30] );
FullAdder eig3fa32( Sev3_C_[31], Sev3_S_[32], Six5_C[25], Eig3_S_[31], Eig3_C_[31] );
FullAdder eig3fa33( Sev3_C_[32], Sev3_S_[33], Six5_C[26], Eig3_S_[32], Eig3_C_[32] );
FullAdder eig3fa34( Sev3_C_[33], Sev3_S_[34], Six5_C[27], Eig3_S_[33], Eig3_C_[33] );
FullAdder eig3fa35( Sev3_C_[34], Six5_S[29], Six5_C[28], Eig3_S_[34], Eig3_C_[34] );
HalfAdder eig3fa36( Six5_S[30], Six5_C[29], Eig3_S_[35], Eig3_C_[35] );
HalfAdder eig3fa37( Six5_S[31], Six5_C[30], Eig3_S_[36], Eig3_C_[36] );

reg	[31: 0]	Eig1_S, Eig1_C;
reg	[35: 0]	Eig2_S, Eig2_C;
reg	[36: 0]	Eig3_S, Eig3_C;

reg done7;
reg state_done7;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Eig1_S <= 32'b0;  Eig1_C <= 32'b0;
    Eig2_S <= 36'b0;  Eig2_C <= 36'b0;
    Eig3_S <= 37'b0;  Eig3_C <= 37'b0;
    done7 <= 1'b0;
    state_done7 <= 1'b0;
  end else begin
    case (state_done7)
      1'b0: begin
        if (done6) begin
          Eig1_S <= Eig1_S_;  Eig1_C <= Eig1_C_;
          Eig2_S <= Eig2_S_;  Eig2_C <= Eig2_C_;
          Eig3_S <= Eig3_S_;  Eig3_C <= Eig3_C_;
          done7 <= 1'b1;
          state_done7 <= 1'b1;
        end else begin
          done7 <= 1'b0;
        end
      end
      1'b1: begin
        done7 <= 1'b0;
        if (!done6)
          state_done7 <= 1'b0;
      end
    endcase
  end
end


//===================Ninth stage===============================

wire	[31: 0]	Nin1_S, Nin1_C;
wire	[41: 0]	Nin2_S, Nin2_C;



HalfAdder nin1fa1( Eig1_C[0], Eig1_S[1], Nin1_S[0], Nin1_C[0] );
HalfAdder nin1fa2( Eig1_C[1], Eig1_S[2], Nin1_S[1], Nin1_C[1] );
HalfAdder nin1fa3( Eig1_C[2], Eig1_S[3], Nin1_S[2], Nin1_C[2] );
HalfAdder nin1fa4( Eig1_C[3], Eig1_S[4], Nin1_S[3], Nin1_C[3] );
FullAdder nin1fa5( Eig1_C[4], Eig1_S[5], Six2_C[0], Nin1_S[4], Nin1_C[4] );
FullAdder nin1fa6( Eig1_C[5], Eig1_S[6], Six2_C[1], Nin1_S[5], Nin1_C[5] );
FullAdder nin1fa7( Eig1_C[6], Eig1_S[7], Six2_C[2], Nin1_S[6], Nin1_C[6] );
FullAdder nin1fa8( Eig1_C[7], Eig1_S[8], Six2_C[3], Nin1_S[7], Nin1_C[7] );
FullAdder nin1fa9(  Eig1_C[8],  Eig1_S[9],  Sev2_S_[0],  Nin1_S[8],  Nin1_C[8] );
FullAdder nin1fa10( Eig1_C[9],  Eig1_S[10], Eig2_S[0],  Nin1_S[9],  Nin1_C[9] );
FullAdder nin1fa11( Eig1_C[10], Eig1_S[11], Eig2_S[1],  Nin1_S[10], Nin1_C[10] );
FullAdder nin1fa12( Eig1_C[11], Eig1_S[12], Eig2_S[2],  Nin1_S[11], Nin1_C[11] );
FullAdder nin1fa13( Eig1_C[12], Eig1_S[13], Eig2_S[3],  Nin1_S[12], Nin1_C[12] );
FullAdder nin1fa14( Eig1_C[13], Eig1_S[14], Eig2_S[4],  Nin1_S[13], Nin1_C[13] );
FullAdder nin1fa15( Eig1_C[14], Eig1_S[15], Eig2_S[5],  Nin1_S[14], Nin1_C[14] );
FullAdder nin1fa16( Eig1_C[15], Eig1_S[16], Eig2_S[6],  Nin1_S[15], Nin1_C[15] );
FullAdder nin1fa17( Eig1_C[16], Eig1_S[17], Eig2_S[7],  Nin1_S[16], Nin1_C[16] );
FullAdder nin1fa18( Eig1_C[17], Eig1_S[18], Eig2_S[8],  Nin1_S[17], Nin1_C[17] );
FullAdder nin1fa19( Eig1_C[18], Eig1_S[19], Eig2_S[9], Nin1_S[18], Nin1_C[18] );
FullAdder nin1fa20( Eig1_C[19], Eig1_S[20], Eig2_S[10], Nin1_S[19], Nin1_C[19] );
FullAdder nin1fa21( Eig1_C[20], Eig1_S[21], Eig2_S[11], Nin1_S[20], Nin1_C[20] );
FullAdder nin1fa22( Eig1_C[21], Eig1_S[22], Eig2_S[12], Nin1_S[21], Nin1_C[21] );
FullAdder nin1fa23( Eig1_C[22], Eig1_S[23], Eig2_S[13], Nin1_S[22], Nin1_C[22] );
FullAdder nin1fa24( Eig1_C[23], Eig1_S[24], Eig2_S[14], Nin1_S[23], Nin1_C[23] );
FullAdder nin1fa25( Eig1_C[24], Eig1_S[25], Eig2_S[15], Nin1_S[24], Nin1_C[24] );
FullAdder nin1fa26( Eig1_C[25], Eig1_S[26], Eig2_S[16], Nin1_S[25], Nin1_C[25] );
FullAdder nin1fa27( Eig1_C[26], Eig1_S[27], Eig2_S[17], Nin1_S[26], Nin1_C[26] );
FullAdder nin1fa28( Eig1_C[27], Eig1_S[28], Eig2_S[18], Nin1_S[27], Nin1_C[27] );
FullAdder nin1fa29( Eig1_C[28], Eig1_S[29], Eig2_S[19], Nin1_S[28], Nin1_C[28] );
FullAdder nin1fa30( Eig1_C[29], Eig1_S[30], Eig2_S[20], Nin1_S[29], Nin1_C[29] );
FullAdder nin1fa31( Eig1_C[30], Eig1_S[31], Eig2_S[21], Nin1_S[30], Nin1_C[30] );
HalfAdder nin1fa32( Eig1_C[31], Eig2_S[22], Nin1_S[31], Nin1_C[31] );


HalfAdder nin2fa1( Eig2_C[6], Fou5_C[0], Nin2_S[0], Nin2_C[0] );
HalfAdder nin2fa2( Eig2_C[7], Fif4_S_[0], Nin2_S[1], Nin2_C[1] );
HalfAdder nin2fa3( Eig2_C[8], Six4_S[0], Nin2_S[2], Nin2_C[2] );
HalfAdder nin2fa4( Eig2_C[9], Sev3_S_[0], Nin2_S[3], Nin2_C[3] );
HalfAdder nin2fa5( Eig2_C[10], Eig3_S[0], Nin2_S[4], Nin2_C[4] );
FullAdder nin2fa6( Eig2_C[11], Eig3_S[1], Eig3_C[0], Nin2_S[5], Nin2_C[5] );
FullAdder nin2fa7( Eig2_C[12], Eig3_S[2], Eig3_C[1], Nin2_S[6], Nin2_C[6] );
FullAdder nin2fa8( Eig2_C[13], Eig3_S[3], Eig3_C[2], Nin2_S[7], Nin2_C[7] );
FullAdder nin2fa9( Eig2_C[14], Eig3_S[4], Eig3_C[3], Nin2_S[8], Nin2_C[8] );
FullAdder nin2fa10( Eig2_C[15], Eig3_S[5], Eig3_C[4], Nin2_S[9], Nin2_C[9] );
FullAdder nin2fa11( Eig2_C[16], Eig3_S[6], Eig3_C[5], Nin2_S[10], Nin2_C[10] );
FullAdder nin2fa12( Eig2_C[17], Eig3_S[7], Eig3_C[6], Nin2_S[11], Nin2_C[11] );
FullAdder nin2fa13( Eig2_C[18], Eig3_S[8], Eig3_C[7], Nin2_S[12], Nin2_C[12] );
FullAdder nin2fa14( Eig2_C[19], Eig3_S[9], Eig3_C[8], Nin2_S[13], Nin2_C[13] );
FullAdder nin2fa15( Eig2_C[20], Eig3_S[10], Eig3_C[9], Nin2_S[14], Nin2_C[14] );
FullAdder nin2fa16( Eig2_C[21], Eig3_S[11], Eig3_C[10], Nin2_S[15], Nin2_C[15] );
FullAdder nin2fa17( Eig2_C[22], Eig3_S[12], Eig3_C[11], Nin2_S[16], Nin2_C[16] );
FullAdder nin2fa18( Eig2_C[23], Eig3_S[13], Eig3_C[12], Nin2_S[17], Nin2_C[17] );
FullAdder nin2fa19( Eig2_C[24], Eig3_S[14], Eig3_C[13], Nin2_S[18], Nin2_C[18] );
FullAdder nin2fa20( Eig2_C[25], Eig3_S[15], Eig3_C[14], Nin2_S[19], Nin2_C[19] );
FullAdder nin2fa21( Eig2_C[26], Eig3_S[16], Eig3_C[15], Nin2_S[20], Nin2_C[20] );
FullAdder nin2fa22( Eig2_C[27], Eig3_S[17], Eig3_C[16], Nin2_S[21], Nin2_C[21] );
FullAdder nin2fa23( Eig2_C[28], Eig3_S[18], Eig3_C[17], Nin2_S[22], Nin2_C[22] );
FullAdder nin2fa24( Eig2_C[29], Eig3_S[19], Eig3_C[18], Nin2_S[23], Nin2_C[23] );
FullAdder nin2fa25( Eig2_C[30], Eig3_S[20], Eig3_C[19], Nin2_S[24], Nin2_C[24] );
FullAdder nin2fa26( Eig2_C[31], Eig3_S[21], Eig3_C[20], Nin2_S[25], Nin2_C[25] );
FullAdder nin2fa27( Eig2_C[32], Eig3_S[22], Eig3_C[21], Nin2_S[26], Nin2_C[26] );
FullAdder nin2fa28( Eig2_C[33], Eig3_S[23], Eig3_C[22], Nin2_S[27], Nin2_C[27] );
FullAdder nin2fa29( Eig2_C[34], Eig3_S[24], Eig3_C[23], Nin2_S[28], Nin2_C[28] );
FullAdder nin2fa30( Eig2_C[35], Eig3_S[25], Eig3_C[24], Nin2_S[29], Nin2_C[29] );
HalfAdder nin2fa31( Eig3_S[26], Eig3_C[25], Nin2_S[30], Nin2_C[30] );
HalfAdder nin2fa32( Eig3_S[27], Eig3_C[26], Nin2_S[31], Nin2_C[31] );
HalfAdder nin2fa33( Eig3_S[28], Eig3_C[27], Nin2_S[32], Nin2_C[32] );
HalfAdder nin2fa34( Eig3_S[29], Eig3_C[28], Nin2_S[33], Nin2_C[33] );
HalfAdder nin2fa35( Eig3_S[30], Eig3_C[29], Nin2_S[34], Nin2_C[34] );
HalfAdder nin2fa36( Eig3_S[31], Eig3_C[30], Nin2_S[35], Nin2_C[35] );
HalfAdder nin2fa37( Eig3_S[32], Eig3_C[31], Nin2_S[36], Nin2_C[36] );
HalfAdder nin2fa38( Eig3_S[33], Eig3_C[32], Nin2_S[37], Nin2_C[37] );
HalfAdder nin2fa39( Eig3_S[34], Eig3_C[33], Nin2_S[38], Nin2_C[38] );
HalfAdder nin2fa40( Eig3_S[35], Eig3_C[34], Nin2_S[39], Nin2_C[39] );
HalfAdder nin2fa41( Eig3_S[36], Eig3_C[35], Nin2_S[40], Nin2_C[40] );
HalfAdder nin2fa42( Six5_C[31], Eig3_C[36], Nin2_S[41], Nin2_C[41] );


reg	[31: 0]	Nin1_S_, Nin1_C_;
reg	[41: 0]	Nin2_S_, Nin2_C_;


reg done8;
reg state_done8;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Nin1_S_ <= 32'b0;  Nin1_C_ <= 32'b0;
    Nin2_S_ <= 42'b0;  Nin2_C_ <= 42'b0;
    done8 <= 1'b0;
    state_done8 <= 1'b0;
  end else begin
    case(state_done8)
      1'b0: begin
        if (done7) begin
          Nin1_S_ <= Nin1_S;  Nin1_C_ <= Nin1_C;
          Nin2_S_ <= Nin2_S;  Nin2_C_ <= Nin2_C;
          done8 <= 1'b1;
          state_done8 <= 1'b1;
        end else
          done8 <= 1'b0;
      end
      1'b1: begin
        done8 <= 1'b0;
        if (!done7)
          state_done8 <= 1'b0;
      end
    endcase
  end
end



//===================Tenth stage===============================



wire	[31: 0]	Ten1_S_, Ten1_C_;
wire	[40: 0]	Ten2_S_, Ten2_C_;

assign Ten1_S_=Nin1_S_;
assign Ten1_C_=Nin1_C_;

HalfAdder ten2fa1( Nin2_S_[1], Nin2_C_[0], Ten2_S_[0], Ten2_C_[0] );
HalfAdder ten2fa2( Nin2_S_[2], Nin2_C_[1], Ten2_S_[1], Ten2_C_[1] );
HalfAdder ten2fa3( Nin2_S_[3], Nin2_C_[2], Ten2_S_[2], Ten2_C_[2] );
HalfAdder ten2fa4( Nin2_S_[4], Nin2_C_[3], Ten2_S_[3], Ten2_C_[3] );
HalfAdder ten2fa5( Nin2_S_[5], Nin2_C_[4], Ten2_S_[4], Ten2_C_[4] );
HalfAdder ten2fa6( Nin2_S_[6], Nin2_C_[5], Ten2_S_[5], Ten2_C_[5] );
HalfAdder ten2fa7( Nin2_S_[7], Nin2_C_[6], Ten2_S_[6], Ten2_C_[6] );
HalfAdder ten2fa8( Nin2_S_[8], Nin2_C_[7], Ten2_S_[7], Ten2_C_[7] );
HalfAdder ten2fa9( Nin2_S_[9], Nin2_C_[8], Ten2_S_[8], Ten2_C_[8] );
HalfAdder ten2fa10( Nin2_S_[10], Nin2_C_[9], Ten2_S_[9], Ten2_C_[9] );
HalfAdder ten2fa11( Nin2_S_[11], Nin2_C_[10], Ten2_S_[10], Ten2_C_[10] );
HalfAdder ten2fa12( Nin2_S_[12], Nin2_C_[11], Ten2_S_[11], Ten2_C_[11] );
HalfAdder ten2fa13( Nin2_S_[13], Nin2_C_[12], Ten2_S_[12], Ten2_C_[12] );
HalfAdder ten2fa14( Nin2_S_[14], Nin2_C_[13], Ten2_S_[13], Ten2_C_[13] );
HalfAdder ten2fa15( Nin2_S_[15], Nin2_C_[14], Ten2_S_[14], Ten2_C_[14] );
FullAdder ten2fa16( Eig2_S[23], Nin2_S_[16], Nin2_C_[15], Ten2_S_[15], Ten2_C_[15] );
FullAdder ten2fa17( Eig2_S[24], Nin2_S_[17], Nin2_C_[16], Ten2_S_[16], Ten2_C_[16] );
FullAdder ten2fa18( Eig2_S[25], Nin2_S_[18], Nin2_C_[17], Ten2_S_[17], Ten2_C_[17] );
FullAdder ten2fa19( Eig2_S[26], Nin2_S_[19], Nin2_C_[18], Ten2_S_[18], Ten2_C_[18] );
FullAdder ten2fa20( Eig2_S[27], Nin2_S_[20], Nin2_C_[19], Ten2_S_[19], Ten2_C_[19] );
FullAdder ten2fa21( Eig2_S[28], Nin2_S_[21], Nin2_C_[20], Ten2_S_[20], Ten2_C_[20] );
FullAdder ten2fa22( Eig2_S[29], Nin2_S_[22], Nin2_C_[21], Ten2_S_[21], Ten2_C_[21] );
FullAdder ten2fa23( Eig2_S[30], Nin2_S_[23], Nin2_C_[22], Ten2_S_[22], Ten2_C_[22] );
FullAdder ten2fa24( Eig2_S[31], Nin2_S_[24], Nin2_C_[23], Ten2_S_[23], Ten2_C_[23] );
FullAdder ten2fa25( Eig2_S[32], Nin2_S_[25], Nin2_C_[24], Ten2_S_[24], Ten2_C_[24] );
FullAdder ten2fa26( Eig2_S[33], Nin2_S_[26], Nin2_C_[25], Ten2_S_[25], Ten2_C_[25] );
FullAdder ten2fa27( Eig2_S[34], Nin2_S_[27], Nin2_C_[26], Ten2_S_[26], Ten2_C_[26] );
FullAdder ten2fa28( Eig2_S[35], Nin2_S_[28], Nin2_C_[27], Ten2_S_[27], Ten2_C_[27] );
HalfAdder ten2fa29( Nin2_S_[29], Nin2_C_[28], Ten2_S_[28], Ten2_C_[28] );
HalfAdder ten2fa30( Nin2_S_[30], Nin2_C_[29], Ten2_S_[29], Ten2_C_[29] );
HalfAdder ten2fa31( Nin2_S_[31], Nin2_C_[30], Ten2_S_[30], Ten2_C_[30] );
HalfAdder ten2fa32( Nin2_S_[32], Nin2_C_[31], Ten2_S_[31], Ten2_C_[31] );
HalfAdder ten2fa33( Nin2_S_[33], Nin2_C_[32], Ten2_S_[32], Ten2_C_[32] );
HalfAdder ten2fa34( Nin2_S_[34], Nin2_C_[33], Ten2_S_[33], Ten2_C_[33] );
HalfAdder ten2fa35( Nin2_S_[35], Nin2_C_[34], Ten2_S_[34], Ten2_C_[34] );
HalfAdder ten2fa36( Nin2_S_[36], Nin2_C_[35], Ten2_S_[35], Ten2_C_[35] );
HalfAdder ten2fa37( Nin2_S_[37], Nin2_C_[36], Ten2_S_[36], Ten2_C_[36] );
HalfAdder ten2fa38( Nin2_S_[38], Nin2_C_[37], Ten2_S_[37], Ten2_C_[37] );
HalfAdder ten2fa39( Nin2_S_[39], Nin2_C_[38], Ten2_S_[38], Ten2_C_[38] );
HalfAdder ten2fa40( Nin2_S_[40], Nin2_C_[39], Ten2_S_[39], Ten2_C_[39] );
HalfAdder ten2fa41( Nin2_S_[41], Nin2_C_[40], Ten2_S_[40], Ten2_C_[40] );


reg	[31: 0]	Ten1_S, Ten1_C;
reg	[40: 0]	Ten2_S, Ten2_C;


reg done9;
reg state_done9;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Ten1_S <= 32'b0;  Ten1_C <= 32'b0;
    Ten2_S <= 41'b0;  Ten2_C <= 41'b0;
    done9 <= 1'b0;
    state_done9 <= 1'b0;
  end else begin
    case (state_done9)
      1'b0: begin
        if (done8) begin
          Ten1_S <= Ten1_S_;  Ten1_C <= Ten1_C_;
          Ten2_S <= Ten2_S_;  Ten2_C <= Ten2_C_;
          done9 <= 1'b1;
          state_done9 <= 1'b1;
        end else begin
          done9 <= 1'b0;
        end
      end
      1'b1: begin
        done9 <= 1'b0;
        if (!done8)
          state_done9 <= 1'b0;
      end
    endcase
  end
end



//===================Eleventh stage===============================

wire	[31: 0]	Ele1_S, Ele1_C;

HalfAdder ele1fa1( Ten1_S[1], Ten1_C[0], Ele1_S[0], Ele1_C[0] );
HalfAdder ele1fa2( Ten1_S[2], Ten1_C[1], Ele1_S[1], Ele1_C[1] );
HalfAdder ele1fa3( Ten1_S[3], Ten1_C[2], Ele1_S[2], Ele1_C[2] );
HalfAdder ele1fa4( Ten1_S[4], Ten1_C[3], Ele1_S[3], Ele1_C[3] );
HalfAdder ele1fa5( Ten1_S[5], Ten1_C[4], Ele1_S[4], Ele1_C[4] );
HalfAdder ele1fa6( Ten1_S[6], Ten1_C[5], Ele1_S[5], Ele1_C[5] );
HalfAdder ele1fa7( Ten1_S[7], Ten1_C[6], Ele1_S[6], Ele1_C[6] );
HalfAdder ele1fa8( Ten1_S[8], Ten1_C[7], Ele1_S[7], Ele1_C[7] );
HalfAdder ele1fa9( Ten1_S[9], Ten1_C[8], Ele1_S[8], Ele1_C[8] );
FullAdder ele1fa10( Ten1_S[10], Ten1_C[9], Eig2_C[0], Ele1_S[9], Ele1_C[9] );
FullAdder ele1fa11( Ten1_S[11], Ten1_C[10], Eig2_C[1], Ele1_S[10], Ele1_C[10] );
FullAdder ele1fa12( Ten1_S[12], Ten1_C[11], Eig2_C[2], Ele1_S[11], Ele1_C[11] );
FullAdder ele1fa13( Ten1_S[13], Ten1_C[12], Eig2_C[3], Ele1_S[12], Ele1_C[12] );
FullAdder ele1fa14( Ten1_S[14], Ten1_C[13], Eig2_C[4], Ele1_S[13], Ele1_C[13] );
FullAdder ele1fa15( Ten1_S[15], Ten1_C[14], Eig2_C[5], Ele1_S[14], Ele1_C[14] );
FullAdder ele1fa16( Ten1_S[16], Ten1_C[15], Nin2_S_[0], Ele1_S[15], Ele1_C[15] );
FullAdder ele1fa17( Ten1_S[17], Ten1_C[16], Ten2_S[0], Ele1_S[16], Ele1_C[16] );
FullAdder ele1fa18( Ten1_S[18], Ten1_C[17], Ten2_S[1], Ele1_S[17], Ele1_C[17] );
FullAdder ele1fa19( Ten1_S[19], Ten1_C[18], Ten2_S[2], Ele1_S[18], Ele1_C[18] );
FullAdder ele1fa20( Ten1_S[20], Ten1_C[19], Ten2_S[3], Ele1_S[19], Ele1_C[19] );
FullAdder ele1fa21( Ten1_S[21], Ten1_C[20], Ten2_S[4], Ele1_S[20], Ele1_C[20] );
FullAdder ele1fa22( Ten1_S[22], Ten1_C[21], Ten2_S[5], Ele1_S[21], Ele1_C[21] );
FullAdder ele1fa23( Ten1_S[23], Ten1_C[22], Ten2_S[6], Ele1_S[22], Ele1_C[22] );
FullAdder ele1fa24( Ten1_S[24], Ten1_C[23], Ten2_S[7], Ele1_S[23], Ele1_C[23] );
FullAdder ele1fa25( Ten1_S[25], Ten1_C[24], Ten2_S[8], Ele1_S[24], Ele1_C[24] );
FullAdder ele1fa26( Ten1_S[26], Ten1_C[25], Ten2_S[9], Ele1_S[25], Ele1_C[25] );
FullAdder ele1fa27( Ten1_S[27], Ten1_C[26], Ten2_S[10], Ele1_S[26], Ele1_C[26] );
FullAdder ele1fa28( Ten1_S[28], Ten1_C[27], Ten2_S[11], Ele1_S[27], Ele1_C[27] );
FullAdder ele1fa29( Ten1_S[29], Ten1_C[28], Ten2_S[12], Ele1_S[28], Ele1_C[28] );
FullAdder ele1fa30( Ten1_S[30], Ten1_C[29], Ten2_S[13], Ele1_S[29], Ele1_C[29] );
FullAdder ele1fa31( Ten1_S[31], Ten1_C[30], Ten2_S[14], Ele1_S[30], Ele1_C[30] );
HalfAdder ele1fa32( Ten1_C[31], Ten2_S[15], Ele1_S[31], Ele1_C[31] );

reg	[31: 0]	Ele1_S_, Ele1_C_;
reg done10;
reg state_done10;

always @(posedge clk or posedge reset) begin
  if (reset) begin
    Ele1_S_ <= 32'b0;  Ele1_C_ <= 32'b0;
    done10 <= 1'b0;
    state_done10 <= 1'b0;
  end else begin
    case(state_done10)
      1'b0: begin
        if (done9) begin
          Ele1_S_ <= Ele1_S;  Ele1_C_ <= Ele1_C;
          done10 <= 1'b1;
          state_done10 <= 1'b1;
        end else
          done10 <= 1'b0;
      end
      1'b1: begin
        done10 <= 1'b0;
        if (!done9)
          state_done10 <= 1'b0;
      end
    endcase
  end
end


//===================Twelfth stage===============================

wire	[56: 0]	Twe1_S_, Twe1_C_;

HalfAdder twe1fa1( Ele1_S_[1], Ele1_C_[0], Twe1_S_[0], Twe1_C_[0] );
HalfAdder twe1fa2( Ele1_S_[2], Ele1_C_[1], Twe1_S_[1], Twe1_C_[1] );
HalfAdder twe1fa3( Ele1_S_[3], Ele1_C_[2], Twe1_S_[2], Twe1_C_[2] );
HalfAdder twe1fa4( Ele1_S_[4], Ele1_C_[3], Twe1_S_[3], Twe1_C_[3] );
HalfAdder twe1fa5( Ele1_S_[5], Ele1_C_[4], Twe1_S_[4], Twe1_C_[4] );
HalfAdder twe1fa6( Ele1_S_[6], Ele1_C_[5], Twe1_S_[5], Twe1_C_[5] );
HalfAdder twe1fa7( Ele1_S_[7], Ele1_C_[6], Twe1_S_[6], Twe1_C_[6] );
HalfAdder twe1fa8( Ele1_S_[8], Ele1_C_[7], Twe1_S_[7], Twe1_C_[7] );
HalfAdder twe1fa9( Ele1_S_[9], Ele1_C_[8], Twe1_S_[8], Twe1_C_[8] );
HalfAdder twe1fa10( Ele1_S_[10], Ele1_C_[9], Twe1_S_[9], Twe1_C_[9] );
HalfAdder twe1fa11( Ele1_S_[11], Ele1_C_[10], Twe1_S_[10], Twe1_C_[10] );
HalfAdder twe1fa12( Ele1_S_[12], Ele1_C_[11], Twe1_S_[11], Twe1_C_[11] );
HalfAdder twe1fa13( Ele1_S_[13], Ele1_C_[12], Twe1_S_[12], Twe1_C_[12] );
HalfAdder twe1fa14( Ele1_S_[14], Ele1_C_[13], Twe1_S_[13], Twe1_C_[13] );
HalfAdder twe1fa15( Ele1_S_[15], Ele1_C_[14], Twe1_S_[14], Twe1_C_[14] );
HalfAdder twe1fa16( Ele1_S_[16], Ele1_C_[15], Twe1_S_[15], Twe1_C_[15] );
FullAdder twe1fa17( Ele1_S_[17], Ele1_C_[16], Ten2_C[0], Twe1_S_[16], Twe1_C_[16] );
FullAdder twe1fa18( Ele1_S_[18], Ele1_C_[17], Ten2_C[1], Twe1_S_[17], Twe1_C_[17] );
FullAdder twe1fa19( Ele1_S_[19], Ele1_C_[18], Ten2_C[2], Twe1_S_[18], Twe1_C_[18] );
FullAdder twe1fa20( Ele1_S_[20], Ele1_C_[19], Ten2_C[3], Twe1_S_[19], Twe1_C_[19] );
FullAdder twe1fa21( Ele1_S_[21], Ele1_C_[20], Ten2_C[4], Twe1_S_[20], Twe1_C_[20] );
FullAdder twe1fa22( Ele1_S_[22], Ele1_C_[21], Ten2_C[5], Twe1_S_[21], Twe1_C_[21] );
FullAdder twe1fa23( Ele1_S_[23], Ele1_C_[22], Ten2_C[6], Twe1_S_[22], Twe1_C_[22] );
FullAdder twe1fa24( Ele1_S_[24], Ele1_C_[23], Ten2_C[7], Twe1_S_[23], Twe1_C_[23] );
FullAdder twe1fa25( Ele1_S_[25], Ele1_C_[24], Ten2_C[8], Twe1_S_[24], Twe1_C_[24] );
FullAdder twe1fa26( Ele1_S_[26], Ele1_C_[25], Ten2_C[9], Twe1_S_[25], Twe1_C_[25] );
FullAdder twe1fa27( Ele1_S_[27], Ele1_C_[26], Ten2_C[10], Twe1_S_[26], Twe1_C_[26] );
FullAdder twe1fa28( Ele1_S_[28], Ele1_C_[27], Ten2_C[11], Twe1_S_[27], Twe1_C_[27] );
FullAdder twe1fa29( Ele1_S_[29], Ele1_C_[28], Ten2_C[12], Twe1_S_[28], Twe1_C_[28] );
FullAdder twe1fa30( Ele1_S_[30], Ele1_C_[29], Ten2_C[13], Twe1_S_[29], Twe1_C_[29] );
FullAdder twe1fa31( Ele1_S_[31], Ele1_C_[30], Ten2_C[14], Twe1_S_[30], Twe1_C_[30] );
FullAdder twe1fa32( Ten2_S[16] , Ele1_C_[31], Ten2_C[15], Twe1_S_[31], Twe1_C_[31] );
HalfAdder twe1fa33( Ten2_S[17], Ten2_C[16], Twe1_S_[32], Twe1_C_[32] );
HalfAdder twe1fa34( Ten2_S[18], Ten2_C[17], Twe1_S_[33], Twe1_C_[33] );
HalfAdder twe1fa35( Ten2_S[19], Ten2_C[18], Twe1_S_[34], Twe1_C_[34] );
HalfAdder twe1fa36( Ten2_S[20], Ten2_C[19], Twe1_S_[35], Twe1_C_[35] );
HalfAdder twe1fa37( Ten2_S[21], Ten2_C[20], Twe1_S_[36], Twe1_C_[36] );
HalfAdder twe1fa38( Ten2_S[22], Ten2_C[21], Twe1_S_[37], Twe1_C_[37] );
HalfAdder twe1fa39( Ten2_S[23], Ten2_C[22], Twe1_S_[38], Twe1_C_[38] );
HalfAdder twe1fa40( Ten2_S[24], Ten2_C[23], Twe1_S_[39], Twe1_C_[39] );
HalfAdder twe1fa41( Ten2_S[25], Ten2_C[24], Twe1_S_[40], Twe1_C_[40] );
HalfAdder twe1fa42( Ten2_S[26], Ten2_C[25], Twe1_S_[41], Twe1_C_[41] );
HalfAdder twe1fa43( Ten2_S[27], Ten2_C[26], Twe1_S_[42], Twe1_C_[42] );
HalfAdder twe1fa44( Ten2_S[28], Ten2_C[27], Twe1_S_[43], Twe1_C_[43] );
HalfAdder twe1fa45( Ten2_S[29], Ten2_C[28], Twe1_S_[44], Twe1_C_[44] );
HalfAdder twe1fa46( Ten2_S[30], Ten2_C[29], Twe1_S_[45], Twe1_C_[45] );
HalfAdder twe1fa47( Ten2_S[31], Ten2_C[30], Twe1_S_[46], Twe1_C_[46] );
HalfAdder twe1fa48( Ten2_S[32], Ten2_C[31], Twe1_S_[47], Twe1_C_[47] );
HalfAdder twe1fa49( Ten2_S[33], Ten2_C[32], Twe1_S_[48], Twe1_C_[48] );
HalfAdder twe1fa50( Ten2_S[34], Ten2_C[33], Twe1_S_[49], Twe1_C_[49] );
HalfAdder twe1fa51( Ten2_S[35], Ten2_C[34], Twe1_S_[50], Twe1_C_[50] );
HalfAdder twe1fa52( Ten2_S[36], Ten2_C[35], Twe1_S_[51], Twe1_C_[51] );
HalfAdder twe1fa53( Ten2_S[37], Ten2_C[36], Twe1_S_[52], Twe1_C_[52] );
HalfAdder twe1fa54( Ten2_S[38], Ten2_C[37], Twe1_S_[53], Twe1_C_[53] );
HalfAdder twe1fa55( Ten2_S[39], Ten2_C[38], Twe1_S_[54], Twe1_C_[54] );
HalfAdder twe1fa56( Ten2_S[40], Ten2_C[39], Twe1_S_[55], Twe1_C_[55] );
HalfAdder twe1fa57( Nin2_C_[41], Ten2_C[40], Twe1_S_[56], Twe1_C_[56] );


always @(posedge clk or posedge reset) begin
    if (reset) begin
        opa <= 64'b0;
        opb <= 64'b0;
        done <= 1'b0;
    end else if (done10) begin
        opa <= { Twe1_S_[54 : 0], Ele1_S_[0], Ten1_S[0], Eig1_S[0],
                 Six1_S[0], Fou1_S[0], Thi1_S_[0], Sec1_S[0], Fir1_S_[0], pp0[0] };
        opb <= { Twe1_C_[53: 0], 10'b0 };
        done <= 1;
    end else begin
        done <= 1'b0;
        opa <= 64'b0;
        opb <= 64'b0;
    end
end




endmodule
